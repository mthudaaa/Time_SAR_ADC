magic
tech sky130A
magscale 1 2
timestamp 1722275450
<< nmos >>
rect -500 -141 500 79
<< ndiff >>
rect -558 67 -500 79
rect -558 -129 -546 67
rect -512 -129 -500 67
rect -558 -141 -500 -129
rect 500 67 558 79
rect 500 -129 512 67
rect 546 -129 558 67
rect 500 -141 558 -129
<< ndiffc >>
rect -546 -129 -512 67
rect 512 -129 546 67
<< poly >>
rect -500 151 500 167
rect -500 117 -484 151
rect 484 117 500 151
rect -500 79 500 117
rect -500 -167 500 -141
<< polycont >>
rect -484 117 484 151
<< locali >>
rect -500 117 -484 151
rect 484 117 500 151
rect -546 67 -512 83
rect -546 -145 -512 -129
rect 512 67 546 83
rect 512 -145 546 -129
<< viali >>
rect -484 117 484 151
rect -546 -129 -512 67
rect 512 -129 546 67
<< metal1 >>
rect -496 151 496 157
rect -496 117 -484 151
rect 484 117 496 151
rect -496 111 496 117
rect -552 67 -506 79
rect -552 -129 -546 67
rect -512 -129 -506 67
rect -552 -141 -506 -129
rect 506 67 552 79
rect 506 -129 512 67
rect 546 -129 552 67
rect 506 -141 552 -129
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.1 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
