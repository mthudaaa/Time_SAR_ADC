magic
tech sky130A
magscale 1 2
timestamp 1723455627
<< viali >>
rect 14013 15045 14047 15079
rect 13737 14977 13771 15011
rect 13599 14909 13633 14943
rect 14105 14909 14139 14943
rect 13461 14773 13495 14807
rect 9965 14569 9999 14603
rect 13921 14569 13955 14603
rect 10701 14501 10735 14535
rect 5641 14365 5675 14399
rect 5917 14365 5951 14399
rect 8953 14365 8987 14399
rect 9229 14365 9263 14399
rect 12909 14365 12943 14399
rect 13185 14365 13219 14399
rect 10977 14297 11011 14331
rect 6653 14229 6687 14263
rect 10517 14229 10551 14263
rect 6009 14025 6043 14059
rect 14105 14025 14139 14059
rect 7573 13957 7607 13991
rect 8585 13957 8619 13991
rect 9321 13957 9355 13991
rect 10140 13957 10174 13991
rect 5273 13889 5307 13923
rect 6469 13889 6503 13923
rect 6653 13889 6687 13923
rect 7389 13889 7423 13923
rect 8033 13889 8067 13923
rect 8401 13889 8435 13923
rect 9137 13889 9171 13923
rect 9873 13889 9907 13923
rect 12265 13889 12299 13923
rect 13369 13889 13403 13923
rect 4997 13821 5031 13855
rect 6745 13821 6779 13855
rect 6929 13821 6963 13855
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 7941 13821 7975 13855
rect 8125 13821 8159 13855
rect 8309 13821 8343 13855
rect 11989 13821 12023 13855
rect 13093 13821 13127 13855
rect 8953 13753 8987 13787
rect 7297 13685 7331 13719
rect 11253 13685 11287 13719
rect 13001 13685 13035 13719
rect 5457 13481 5491 13515
rect 5917 13481 5951 13515
rect 8217 13481 8251 13515
rect 8677 13481 8711 13515
rect 12449 13481 12483 13515
rect 13277 13481 13311 13515
rect 6009 13413 6043 13447
rect 6469 13413 6503 13447
rect 6561 13413 6595 13447
rect 8125 13413 8159 13447
rect 8309 13413 8343 13447
rect 10609 13413 10643 13447
rect 9781 13345 9815 13379
rect 10701 13345 10735 13379
rect 12613 13345 12647 13379
rect 13829 13345 13863 13379
rect 5733 13277 5767 13311
rect 5825 13277 5859 13311
rect 6193 13277 6227 13311
rect 6377 13277 6411 13311
rect 6653 13277 6687 13311
rect 6745 13277 6779 13311
rect 7205 13277 7239 13311
rect 7573 13277 7607 13311
rect 7941 13277 7975 13311
rect 8401 13277 8435 13311
rect 9965 13277 9999 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 10977 13277 11011 13311
rect 11253 13277 11287 13311
rect 11345 13277 11379 13311
rect 12725 13277 12759 13311
rect 13415 13277 13449 13311
rect 13553 13277 13587 13311
rect 7389 13209 7423 13243
rect 13001 13209 13035 13243
rect 13093 13209 13127 13243
rect 13921 13209 13955 13243
rect 7021 13141 7055 13175
rect 11253 13141 11287 13175
rect 6469 12869 6503 12903
rect 7021 12869 7055 12903
rect 7113 12869 7147 12903
rect 6653 12801 6687 12835
rect 6745 12733 6779 12767
rect 6929 12733 6963 12767
rect 6469 12393 6503 12427
rect 7941 12393 7975 12427
rect 13461 12393 13495 12427
rect 13829 12257 13863 12291
rect 6377 12189 6411 12223
rect 7849 12189 7883 12223
rect 13645 12189 13679 12223
rect 13921 12189 13955 12223
rect 6469 11101 6503 11135
rect 9965 11101 9999 11135
rect 10241 11101 10275 11135
rect 12541 11101 12575 11135
rect 12817 11101 12851 11135
rect 6285 11033 6319 11067
rect 6653 11033 6687 11067
rect 10977 10965 11011 10999
rect 13553 10965 13587 10999
rect 5917 10761 5951 10795
rect 14013 10761 14047 10795
rect 7573 10693 7607 10727
rect 10609 10693 10643 10727
rect 11069 10693 11103 10727
rect 14565 10693 14599 10727
rect 4905 10625 4939 10659
rect 5181 10625 5215 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7665 10625 7699 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8677 10625 8711 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 10793 10625 10827 10659
rect 10977 10625 11011 10659
rect 13093 10625 13127 10659
rect 14289 10625 14323 10659
rect 7021 10557 7055 10591
rect 7757 10557 7791 10591
rect 7941 10557 7975 10591
rect 8401 10557 8435 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 10241 10557 10275 10591
rect 12817 10557 12851 10591
rect 14177 10557 14211 10591
rect 14657 10557 14691 10591
rect 9781 10489 9815 10523
rect 13829 10489 13863 10523
rect 6469 10421 6503 10455
rect 6837 10421 6871 10455
rect 9413 10421 9447 10455
rect 5733 10217 5767 10251
rect 7021 10217 7055 10251
rect 9045 10217 9079 10251
rect 12909 10217 12943 10251
rect 10057 10149 10091 10183
rect 6193 10081 6227 10115
rect 6837 10081 6871 10115
rect 9413 10081 9447 10115
rect 9505 10081 9539 10115
rect 13461 10081 13495 10115
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 6377 10013 6411 10047
rect 6745 10013 6779 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9689 10013 9723 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 13073 10013 13107 10047
rect 13185 10013 13219 10047
rect 7113 9945 7147 9979
rect 13553 9945 13587 9979
rect 6561 9877 6595 9911
rect 6929 9673 6963 9707
rect 7021 9673 7055 9707
rect 6561 9605 6595 9639
rect 7113 9537 7147 9571
rect 6820 9469 6854 9503
rect 6377 9333 6411 9367
rect 6837 9129 6871 9163
rect 6653 8993 6687 9027
rect 10149 8993 10183 9027
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 6009 8925 6043 8959
rect 6285 8925 6319 8959
rect 10425 8925 10459 8959
rect 12909 8925 12943 8959
rect 13185 8925 13219 8959
rect 6929 8857 6963 8891
rect 7113 8857 7147 8891
rect 5457 8789 5491 8823
rect 11161 8789 11195 8823
rect 13921 8789 13955 8823
rect 10425 8585 10459 8619
rect 11713 8585 11747 8619
rect 13461 8585 13495 8619
rect 12265 8517 12299 8551
rect 14013 8517 14047 8551
rect 10609 8449 10643 8483
rect 10701 8449 10735 8483
rect 10885 8449 10919 8483
rect 10977 8449 11011 8483
rect 11713 8449 11747 8483
rect 13737 8449 13771 8483
rect 11621 8381 11655 8415
rect 13599 8381 13633 8415
rect 14105 8381 14139 8415
rect 7849 8041 7883 8075
rect 7757 7837 7791 7871
rect 8309 7497 8343 7531
rect 12541 7497 12575 7531
rect 6653 7429 6687 7463
rect 8125 7429 8159 7463
rect 11253 7429 11287 7463
rect 6837 7361 6871 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 11345 7361 11379 7395
rect 11805 7361 11839 7395
rect 13533 7361 13567 7395
rect 13645 7361 13679 7395
rect 11529 7293 11563 7327
rect 13921 7293 13955 7327
rect 14013 7293 14047 7327
rect 7021 7225 7055 7259
rect 7389 7157 7423 7191
rect 8309 7157 8343 7191
rect 8493 7157 8527 7191
rect 13369 7157 13403 7191
rect 6193 6953 6227 6987
rect 8401 6953 8435 6987
rect 11437 6953 11471 6987
rect 6728 6817 6762 6851
rect 9413 6817 9447 6851
rect 9505 6817 9539 6851
rect 11069 6817 11103 6851
rect 12587 6817 12621 6851
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 6285 6749 6319 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 9229 6749 9263 6783
rect 9321 6749 9355 6783
rect 9689 6749 9723 6783
rect 10023 6749 10057 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 12449 6749 12483 6783
rect 12909 6749 12943 6783
rect 13185 6719 13219 6753
rect 6469 6681 6503 6715
rect 9781 6681 9815 6715
rect 12081 6681 12115 6715
rect 12173 6681 12207 6715
rect 6837 6613 6871 6647
rect 9045 6613 9079 6647
rect 10609 6613 10643 6647
rect 12725 6613 12759 6647
rect 13921 6613 13955 6647
rect 6193 6409 6227 6443
rect 6837 6409 6871 6443
rect 7757 6409 7791 6443
rect 10609 6409 10643 6443
rect 5181 6273 5215 6307
rect 5457 6273 5491 6307
rect 6745 6273 6779 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 7849 6273 7883 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 13369 6273 13403 6307
rect 6929 6205 6963 6239
rect 13093 6205 13127 6239
rect 6377 6137 6411 6171
rect 14105 6137 14139 6171
rect 10701 5321 10735 5355
rect 11161 5321 11195 5355
rect 10609 5253 10643 5287
rect 10793 5185 10827 5219
rect 11345 5117 11379 5151
rect 11345 4777 11379 4811
rect 11529 4709 11563 4743
rect 10885 4641 10919 4675
rect 9781 4573 9815 4607
rect 10057 4573 10091 4607
rect 10977 4573 11011 4607
rect 11345 4573 11379 4607
rect 9689 4505 9723 4539
rect 9220 4233 9254 4267
rect 8677 4097 8711 4131
rect 8861 4097 8895 4131
rect 9597 4097 9631 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 10701 4097 10735 4131
rect 10793 4097 10827 4131
rect 13553 4097 13587 4131
rect 13829 4097 13863 4131
rect 10149 4029 10183 4063
rect 12817 4029 12851 4063
rect 13461 4029 13495 4063
rect 8585 3961 8619 3995
rect 9781 3961 9815 3995
rect 13185 3961 13219 3995
rect 9045 3893 9079 3927
rect 9229 3893 9263 3927
rect 13277 3893 13311 3927
rect 8677 3689 8711 3723
rect 10701 3689 10735 3723
rect 13829 3689 13863 3723
rect 14197 3689 14231 3723
rect 12265 3553 12299 3587
rect 12449 3553 12483 3587
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 9338 3485 9372 3519
rect 9597 3485 9631 3519
rect 9689 3485 9723 3519
rect 9965 3485 9999 3519
rect 12357 3485 12391 3519
rect 12716 3485 12750 3519
rect 14289 3485 14323 3519
rect 14381 3145 14415 3179
rect 13268 3077 13302 3111
rect 8861 3009 8895 3043
rect 9137 3009 9171 3043
rect 13001 2941 13035 2975
rect 9873 2805 9907 2839
<< metal1 >>
rect 1104 15802 15088 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 15088 15802
rect 1104 15728 15088 15750
rect 1104 15258 15088 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 15088 15258
rect 1104 15184 15088 15206
rect 13998 15036 14004 15088
rect 14056 15036 14062 15088
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 13587 14943 13645 14949
rect 13587 14940 13599 14943
rect 12216 14912 13599 14940
rect 12216 14900 12222 14912
rect 13587 14909 13599 14912
rect 13633 14909 13645 14943
rect 13587 14903 13645 14909
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 13078 14832 13084 14884
rect 13136 14872 13142 14884
rect 14108 14872 14136 14903
rect 13136 14844 14136 14872
rect 13136 14832 13142 14844
rect 13170 14764 13176 14816
rect 13228 14804 13234 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 13228 14776 13461 14804
rect 13228 14764 13234 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 13449 14767 13507 14773
rect 1104 14714 15088 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 15088 14714
rect 1104 14640 15088 14662
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9364 14572 9965 14600
rect 9364 14560 9370 14572
rect 9953 14569 9965 14572
rect 9999 14600 10011 14603
rect 12158 14600 12164 14612
rect 9999 14572 12164 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 13909 14603 13967 14609
rect 13909 14569 13921 14603
rect 13955 14600 13967 14603
rect 13998 14600 14004 14612
rect 13955 14572 14004 14600
rect 13955 14569 13967 14572
rect 13909 14563 13967 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 10686 14492 10692 14544
rect 10744 14532 10750 14544
rect 11054 14532 11060 14544
rect 10744 14504 11060 14532
rect 10744 14492 10750 14504
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 4672 14368 5641 14396
rect 4672 14356 4678 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5644 14328 5672 14359
rect 5902 14356 5908 14408
rect 5960 14356 5966 14408
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 8956 14328 8984 14359
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13078 14396 13084 14408
rect 12943 14368 13084 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13170 14356 13176 14408
rect 13228 14356 13234 14408
rect 9766 14328 9772 14340
rect 5644 14300 9772 14328
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 10870 14288 10876 14340
rect 10928 14328 10934 14340
rect 10965 14331 11023 14337
rect 10965 14328 10977 14331
rect 10928 14300 10977 14328
rect 10928 14288 10934 14300
rect 10965 14297 10977 14300
rect 11011 14297 11023 14331
rect 10965 14291 11023 14297
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 7558 14260 7564 14272
rect 6687 14232 7564 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 1104 14170 15088 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 15088 14170
rect 1104 14096 15088 14118
rect 5997 14059 6055 14065
rect 5997 14025 6009 14059
rect 6043 14056 6055 14059
rect 12618 14056 12624 14068
rect 6043 14028 12624 14056
rect 6043 14025 6055 14028
rect 5997 14019 6055 14025
rect 5442 13948 5448 14000
rect 5500 13988 5506 14000
rect 7576 13997 7604 14028
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 7561 13991 7619 13997
rect 5500 13960 6684 13988
rect 5500 13948 5506 13960
rect 6656 13929 6684 13960
rect 6932 13960 7512 13988
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 5307 13892 6469 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 6457 13883 6515 13889
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6932 13920 6960 13960
rect 6641 13883 6699 13889
rect 6840 13892 6960 13920
rect 4614 13812 4620 13864
rect 4672 13852 4678 13864
rect 4985 13855 5043 13861
rect 4985 13852 4997 13855
rect 4672 13824 4997 13852
rect 4672 13812 4678 13824
rect 4985 13821 4997 13824
rect 5031 13821 5043 13855
rect 4985 13815 5043 13821
rect 6730 13812 6736 13864
rect 6788 13812 6794 13864
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 6840 13784 6868 13892
rect 7374 13880 7380 13932
rect 7432 13880 7438 13932
rect 7484 13920 7512 13960
rect 7561 13957 7573 13991
rect 7607 13957 7619 13991
rect 7561 13951 7619 13957
rect 8573 13991 8631 13997
rect 8573 13957 8585 13991
rect 8619 13988 8631 13991
rect 9214 13988 9220 14000
rect 8619 13960 9220 13988
rect 8619 13957 8631 13960
rect 8573 13951 8631 13957
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 9306 13948 9312 14000
rect 9364 13948 9370 14000
rect 10128 13991 10186 13997
rect 10128 13957 10140 13991
rect 10174 13988 10186 13991
rect 13446 13988 13452 14000
rect 10174 13960 13452 13988
rect 10174 13957 10186 13960
rect 10128 13951 10186 13957
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 7650 13920 7656 13932
rect 7484 13892 7656 13920
rect 7650 13880 7656 13892
rect 7708 13920 7714 13932
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 7708 13892 8033 13920
rect 7708 13880 7714 13892
rect 8021 13889 8033 13892
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 8662 13920 8668 13932
rect 8435 13892 8668 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 9048 13892 9137 13920
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7834 13852 7840 13864
rect 7147 13824 7840 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 7926 13812 7932 13864
rect 7984 13812 7990 13864
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8478 13852 8484 13864
rect 8343 13824 8484 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8128 13784 8156 13815
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 6512 13756 6868 13784
rect 7116 13756 8156 13784
rect 6512 13744 6518 13756
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7116 13716 7144 13756
rect 8386 13744 8392 13796
rect 8444 13784 8450 13796
rect 8941 13787 8999 13793
rect 8941 13784 8953 13787
rect 8444 13756 8953 13784
rect 8444 13744 8450 13756
rect 8941 13753 8953 13756
rect 8987 13753 8999 13787
rect 8941 13747 8999 13753
rect 6972 13688 7144 13716
rect 6972 13676 6978 13688
rect 7282 13676 7288 13728
rect 7340 13676 7346 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 9048 13716 9076 13892
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10502 13920 10508 13932
rect 9907 13892 10508 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12434 13920 12440 13932
rect 12299 13892 12440 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 10226 13716 10232 13728
rect 7524 13688 10232 13716
rect 7524 13676 7530 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 11238 13676 11244 13728
rect 11296 13676 11302 13728
rect 11992 13716 12020 13815
rect 13078 13812 13084 13864
rect 13136 13812 13142 13864
rect 13096 13784 13124 13812
rect 12544 13756 13124 13784
rect 12544 13716 12572 13756
rect 11992 13688 12572 13716
rect 12986 13676 12992 13728
rect 13044 13676 13050 13728
rect 1104 13626 15088 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 15088 13626
rect 1104 13552 15088 13574
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 5905 13515 5963 13521
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 6822 13512 6828 13524
rect 5951 13484 6828 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 6822 13472 6828 13484
rect 6880 13512 6886 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 6880 13484 8217 13512
rect 6880 13472 6886 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8205 13475 8263 13481
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 13265 13515 13323 13521
rect 13265 13481 13277 13515
rect 13311 13512 13323 13515
rect 13354 13512 13360 13524
rect 13311 13484 13360 13512
rect 13311 13481 13323 13484
rect 13265 13475 13323 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 5997 13447 6055 13453
rect 5997 13413 6009 13447
rect 6043 13444 6055 13447
rect 6454 13444 6460 13456
rect 6043 13416 6460 13444
rect 6043 13413 6055 13416
rect 5997 13407 6055 13413
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 6549 13447 6607 13453
rect 6549 13413 6561 13447
rect 6595 13444 6607 13447
rect 6914 13444 6920 13456
rect 6595 13416 6920 13444
rect 6595 13413 6607 13416
rect 6549 13407 6607 13413
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 7064 13416 8125 13444
rect 7064 13404 7070 13416
rect 8113 13413 8125 13416
rect 8159 13413 8171 13447
rect 8113 13407 8171 13413
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13444 8355 13447
rect 10597 13447 10655 13453
rect 10597 13444 10609 13447
rect 8343 13416 10609 13444
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 10597 13413 10609 13416
rect 10643 13413 10655 13447
rect 10597 13407 10655 13413
rect 7282 13376 7288 13388
rect 5736 13348 7288 13376
rect 5736 13317 5764 13348
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 8018 13336 8024 13388
rect 8076 13376 8082 13388
rect 8312 13376 8340 13407
rect 8076 13348 8340 13376
rect 8076 13336 8082 13348
rect 9766 13336 9772 13388
rect 9824 13336 9830 13388
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 10152 13348 10701 13376
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13308 6239 13311
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6227 13280 6377 13308
rect 6227 13277 6239 13280
rect 6181 13271 6239 13277
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 5828 13172 5856 13271
rect 6380 13240 6408 13271
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 6604 13280 6653 13308
rect 6604 13268 6610 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6779 13280 7205 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 7558 13268 7564 13320
rect 7616 13268 7622 13320
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7892 13280 7941 13308
rect 7892 13268 7898 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 10152 13317 10180 13348
rect 10689 13345 10701 13348
rect 10735 13376 10747 13379
rect 10870 13376 10876 13388
rect 10735 13348 10876 13376
rect 10735 13345 10747 13348
rect 10689 13339 10747 13345
rect 10870 13336 10876 13348
rect 10928 13376 10934 13388
rect 11698 13376 11704 13388
rect 10928 13348 11704 13376
rect 10928 13336 10934 13348
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12618 13385 12624 13388
rect 12601 13379 12624 13385
rect 12601 13345 12613 13379
rect 12601 13339 12624 13345
rect 12618 13336 12624 13339
rect 12676 13336 12682 13388
rect 13817 13379 13875 13385
rect 12728 13348 13584 13376
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 8536 13280 9965 13308
rect 8536 13268 8542 13280
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 7377 13243 7435 13249
rect 6380 13212 7144 13240
rect 6546 13172 6552 13184
rect 5828 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6696 13144 7021 13172
rect 6696 13132 6702 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7116 13172 7144 13212
rect 7377 13209 7389 13243
rect 7423 13240 7435 13243
rect 7466 13240 7472 13252
rect 7423 13212 7472 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 7926 13172 7932 13184
rect 7116 13144 7932 13172
rect 7009 13135 7067 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9968 13172 9996 13271
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 10284 13280 10333 13308
rect 10284 13268 10290 13280
rect 10321 13277 10333 13280
rect 10367 13308 10379 13311
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10367 13280 10977 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 12728 13317 12756 13348
rect 13556 13317 13584 13348
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 14090 13376 14096 13388
rect 13863 13348 14096 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13277 12771 13311
rect 13403 13311 13461 13317
rect 13403 13308 13415 13311
rect 12713 13271 12771 13277
rect 12820 13280 13415 13308
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11348 13240 11376 13271
rect 11204 13212 11376 13240
rect 11204 13200 11210 13212
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 12250 13240 12256 13252
rect 11480 13212 12256 13240
rect 11480 13200 11486 13212
rect 12250 13200 12256 13212
rect 12308 13240 12314 13252
rect 12820 13240 12848 13280
rect 13403 13277 13415 13280
rect 13449 13277 13461 13311
rect 13403 13271 13461 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 13722 13308 13728 13320
rect 13587 13280 13728 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 12308 13212 12848 13240
rect 12308 13200 12314 13212
rect 12986 13200 12992 13252
rect 13044 13200 13050 13252
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 13909 13243 13967 13249
rect 13909 13240 13921 13243
rect 13136 13212 13921 13240
rect 13136 13200 13142 13212
rect 13909 13209 13921 13212
rect 13955 13209 13967 13243
rect 13909 13203 13967 13209
rect 11238 13172 11244 13184
rect 9968 13144 11244 13172
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 13096 13172 13124 13200
rect 12768 13144 13124 13172
rect 12768 13132 12774 13144
rect 1104 13082 15088 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 15088 13082
rect 1104 13008 15088 13030
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 8018 12968 8024 12980
rect 6604 12940 8024 12968
rect 6604 12928 6610 12940
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 5902 12860 5908 12912
rect 5960 12900 5966 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 5960 12872 6469 12900
rect 5960 12860 5966 12872
rect 6457 12869 6469 12872
rect 6503 12869 6515 12903
rect 6457 12863 6515 12869
rect 7006 12860 7012 12912
rect 7064 12860 7070 12912
rect 7101 12903 7159 12909
rect 7101 12869 7113 12903
rect 7147 12900 7159 12903
rect 7834 12900 7840 12912
rect 7147 12872 7840 12900
rect 7147 12869 7159 12872
rect 7101 12863 7159 12869
rect 7834 12860 7840 12872
rect 7892 12860 7898 12912
rect 6638 12792 6644 12844
rect 6696 12792 6702 12844
rect 7024 12832 7052 12860
rect 7374 12832 7380 12844
rect 7024 12804 7380 12832
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 11422 12832 11428 12844
rect 7616 12804 11428 12832
rect 7616 12792 7622 12804
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 6730 12724 6736 12776
rect 6788 12724 6794 12776
rect 6822 12724 6828 12776
rect 6880 12764 6886 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6880 12736 6929 12764
rect 6880 12724 6886 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 6748 12696 6776 12724
rect 8478 12696 8484 12708
rect 6748 12668 8484 12696
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 1104 12538 15088 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 15088 12538
rect 1104 12464 15088 12486
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 6822 12424 6828 12436
rect 6503 12396 6828 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7926 12384 7932 12436
rect 7984 12384 7990 12436
rect 13446 12384 13452 12436
rect 13504 12384 13510 12436
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12288 13875 12291
rect 14182 12288 14188 12300
rect 13863 12260 14188 12288
rect 13863 12257 13875 12260
rect 13817 12251 13875 12257
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6914 12220 6920 12232
rect 6411 12192 6920 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 10318 12180 10324 12232
rect 10376 12220 10382 12232
rect 13633 12223 13691 12229
rect 13633 12220 13645 12223
rect 10376 12192 13645 12220
rect 10376 12180 10382 12192
rect 13633 12189 13645 12192
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 13648 12152 13676 12183
rect 13906 12180 13912 12232
rect 13964 12180 13970 12232
rect 13814 12152 13820 12164
rect 13648 12124 13820 12152
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 1104 11994 15088 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 15088 11994
rect 1104 11920 15088 11942
rect 1104 11450 15088 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 15088 11450
rect 1104 11376 15088 11398
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 7466 11132 7472 11144
rect 6503 11104 7472 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9824 11104 9965 11132
rect 9824 11092 9830 11104
rect 9953 11101 9965 11104
rect 9999 11132 10011 11135
rect 10134 11132 10140 11144
rect 9999 11104 10140 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12710 11132 12716 11144
rect 12575 11104 12716 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12802 11092 12808 11144
rect 12860 11092 12866 11144
rect 6273 11067 6331 11073
rect 6273 11033 6285 11067
rect 6319 11033 6331 11067
rect 6273 11027 6331 11033
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 6730 11064 6736 11076
rect 6687 11036 6736 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6288 10996 6316 11027
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 10888 11036 11100 11064
rect 10888 10996 10916 11036
rect 5960 10968 10916 10996
rect 5960 10956 5966 10968
rect 10962 10956 10968 11008
rect 11020 10956 11026 11008
rect 11072 10996 11100 11036
rect 12342 10996 12348 11008
rect 11072 10968 12348 10996
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 13538 10956 13544 11008
rect 13596 10956 13602 11008
rect 1104 10906 15088 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 15088 10906
rect 1104 10832 15088 10854
rect 5902 10752 5908 10804
rect 5960 10752 5966 10804
rect 7006 10792 7012 10804
rect 6656 10764 7012 10792
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4672 10628 4905 10656
rect 4672 10616 4678 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5718 10656 5724 10668
rect 5215 10628 5724 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6144 10424 6469 10452
rect 6144 10412 6150 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6656 10452 6684 10764
rect 7006 10752 7012 10764
rect 7064 10792 7070 10804
rect 8018 10792 8024 10804
rect 7064 10764 8024 10792
rect 7064 10752 7070 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 10962 10752 10968 10804
rect 11020 10752 11026 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13096 10764 14013 10792
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 7926 10724 7932 10736
rect 7607 10696 7932 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7576 10656 7604 10687
rect 7926 10684 7932 10696
rect 7984 10684 7990 10736
rect 8036 10724 8064 10752
rect 8036 10696 10180 10724
rect 7239 10628 7604 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7650 10616 7656 10668
rect 7708 10616 7714 10668
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 10152 10665 10180 10696
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10597 10727 10655 10733
rect 10597 10724 10609 10727
rect 10284 10696 10609 10724
rect 10284 10684 10290 10696
rect 10597 10693 10609 10696
rect 10643 10693 10655 10727
rect 10980 10724 11008 10752
rect 10597 10687 10655 10693
rect 10704 10696 11008 10724
rect 11057 10727 11115 10733
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8251 10628 8677 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10704 10656 10732 10696
rect 11057 10693 11069 10727
rect 11103 10724 11115 10727
rect 11238 10724 11244 10736
rect 11103 10696 11244 10724
rect 11103 10693 11115 10696
rect 11057 10687 11115 10693
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 10459 10628 10732 10656
rect 10781 10659 10839 10665
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 6822 10548 6828 10600
rect 6880 10548 6886 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7374 10588 7380 10600
rect 7055 10560 7380 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 6840 10520 6868 10548
rect 7760 10520 7788 10551
rect 7926 10548 7932 10600
rect 7984 10548 7990 10600
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 9858 10588 9864 10600
rect 9324 10560 9864 10588
rect 6840 10492 7788 10520
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6656 10424 6837 10452
rect 6457 10415 6515 10421
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 9324 10452 9352 10560
rect 9858 10548 9864 10560
rect 9916 10588 9922 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9916 10560 9965 10588
rect 9916 10548 9922 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 10796 10520 10824 10619
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 13096 10665 13124 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 13780 10696 14320 10724
rect 13780 10684 13786 10696
rect 14292 10665 14320 10696
rect 14550 10684 14556 10736
rect 14608 10684 14614 10736
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10928 10628 10977 10656
rect 10928 10616 10934 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12768 10560 12817 10588
rect 12768 10548 12774 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 14165 10591 14223 10597
rect 14165 10588 14177 10591
rect 12805 10551 12863 10557
rect 13464 10560 14177 10588
rect 9815 10492 10824 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 7708 10424 9352 10452
rect 9401 10455 9459 10461
rect 7708 10412 7714 10424
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 9490 10452 9496 10464
rect 9447 10424 9496 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 9490 10412 9496 10424
rect 9548 10452 9554 10464
rect 13464 10452 13492 10560
rect 14165 10557 14177 10560
rect 14211 10588 14223 10591
rect 14366 10588 14372 10600
rect 14211 10560 14372 10588
rect 14211 10557 14223 10560
rect 14165 10551 14223 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 13817 10523 13875 10529
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 14550 10520 14556 10532
rect 13863 10492 14556 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 14550 10480 14556 10492
rect 14608 10480 14614 10532
rect 9548 10424 13492 10452
rect 9548 10412 9554 10424
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14660 10452 14688 10551
rect 14148 10424 14688 10452
rect 14148 10412 14154 10424
rect 1104 10362 15088 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 15088 10362
rect 1104 10288 15088 10310
rect 5718 10208 5724 10260
rect 5776 10208 5782 10260
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6328 10220 7021 10248
rect 6328 10208 6334 10220
rect 7009 10217 7021 10220
rect 7055 10248 7067 10251
rect 7650 10248 7656 10260
rect 7055 10220 7656 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 8076 10220 9045 10248
rect 8076 10208 8082 10220
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 9033 10211 9091 10217
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12860 10220 12909 10248
rect 12860 10208 12866 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 12897 10211 12955 10217
rect 4614 10140 4620 10192
rect 4672 10180 4678 10192
rect 8386 10180 8392 10192
rect 4672 10152 8392 10180
rect 4672 10140 4678 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 10045 10183 10103 10189
rect 10045 10149 10057 10183
rect 10091 10180 10103 10183
rect 10870 10180 10876 10192
rect 10091 10152 10876 10180
rect 10091 10149 10103 10152
rect 10045 10143 10103 10149
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 6086 10112 6092 10124
rect 5920 10084 6092 10112
rect 5920 10053 5948 10084
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6822 10112 6828 10124
rect 6227 10084 6828 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6822 10072 6828 10084
rect 6880 10112 6886 10124
rect 6880 10084 7236 10112
rect 6880 10072 6886 10084
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 5994 10004 6000 10056
rect 6052 10004 6058 10056
rect 6270 10004 6276 10056
rect 6328 10004 6334 10056
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6411 10016 6745 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 6733 10013 6745 10016
rect 6779 10044 6791 10047
rect 6779 10016 6960 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 6546 9868 6552 9920
rect 6604 9868 6610 9920
rect 6932 9908 6960 10016
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7208 10053 7236 10084
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 7432 10084 7972 10112
rect 7432 10072 7438 10084
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7834 10044 7840 10056
rect 7515 10016 7840 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 7190 9908 7196 9920
rect 6932 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9908 7254 9920
rect 7484 9908 7512 10007
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 7944 10044 7972 10084
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 9401 10115 9459 10121
rect 9401 10112 9413 10115
rect 8168 10084 9413 10112
rect 8168 10072 8174 10084
rect 9401 10081 9413 10084
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 9490 10072 9496 10124
rect 9548 10072 9554 10124
rect 10226 10112 10232 10124
rect 9692 10084 10232 10112
rect 9692 10056 9720 10084
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 7944 10016 9229 10044
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 7558 9936 7564 9988
rect 7616 9976 7622 9988
rect 9324 9976 9352 10007
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 10042 10004 10048 10056
rect 10100 10004 10106 10056
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 13078 10053 13084 10056
rect 13061 10047 13084 10053
rect 13061 10044 13073 10047
rect 11020 10016 13073 10044
rect 11020 10004 11026 10016
rect 13061 10013 13073 10016
rect 13061 10007 13084 10013
rect 13078 10004 13084 10007
rect 13136 10004 13142 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13722 10044 13728 10056
rect 13219 10016 13728 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 10060 9976 10088 10004
rect 7616 9948 10088 9976
rect 7616 9936 7622 9948
rect 12710 9936 12716 9988
rect 12768 9976 12774 9988
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 12768 9948 13553 9976
rect 12768 9936 12774 9948
rect 13541 9945 13553 9948
rect 13587 9976 13599 9979
rect 14090 9976 14096 9988
rect 13587 9948 14096 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 7248 9880 7512 9908
rect 7248 9868 7254 9880
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 11238 9908 11244 9920
rect 7984 9880 11244 9908
rect 7984 9868 7990 9880
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 1104 9818 15088 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 15088 9818
rect 1104 9744 15088 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6052 9676 6868 9704
rect 6052 9664 6058 9676
rect 6546 9596 6552 9648
rect 6604 9596 6610 9648
rect 6840 9636 6868 9676
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 7009 9707 7067 9713
rect 7009 9673 7021 9707
rect 7055 9704 7067 9707
rect 7926 9704 7932 9716
rect 7055 9676 7932 9704
rect 7055 9673 7067 9676
rect 7009 9667 7067 9673
rect 7024 9636 7052 9667
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 6840 9608 7052 9636
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 9674 9636 9680 9648
rect 7524 9608 9680 9636
rect 7524 9596 7530 9608
rect 9674 9596 9680 9608
rect 9732 9636 9738 9648
rect 10962 9636 10968 9648
rect 9732 9608 10968 9636
rect 9732 9596 9738 9608
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 6822 9509 6828 9512
rect 6808 9503 6828 9509
rect 6808 9469 6820 9503
rect 6808 9463 6828 9469
rect 6822 9460 6828 9463
rect 6880 9460 6886 9512
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 4764 9336 6377 9364
rect 4764 9324 4770 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 1104 9274 15088 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 15088 9274
rect 1104 9200 15088 9222
rect 6822 9120 6828 9172
rect 6880 9120 6886 9172
rect 7374 9092 7380 9104
rect 6012 9064 7380 9092
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 4614 8956 4620 8968
rect 4479 8928 4620 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 6012 8965 6040 9064
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 6914 9024 6920 9036
rect 6687 8996 6920 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 10134 8984 10140 9036
rect 10192 8984 10198 9036
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8956 6331 8959
rect 7558 8956 7564 8968
rect 6319 8928 7564 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 6914 8848 6920 8900
rect 6972 8848 6978 8900
rect 7101 8891 7159 8897
rect 7101 8857 7113 8891
rect 7147 8888 7159 8891
rect 12618 8888 12624 8900
rect 7147 8860 12624 8888
rect 7147 8857 7159 8860
rect 7101 8851 7159 8857
rect 5445 8823 5503 8829
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 7116 8820 7144 8851
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 12912 8888 12940 8919
rect 13170 8916 13176 8968
rect 13228 8916 13234 8968
rect 14090 8888 14096 8900
rect 12912 8860 14096 8888
rect 14090 8848 14096 8860
rect 14148 8848 14154 8900
rect 5491 8792 7144 8820
rect 11149 8823 11207 8829
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 12434 8820 12440 8832
rect 11195 8792 12440 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13906 8780 13912 8832
rect 13964 8780 13970 8832
rect 1104 8730 15088 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 15088 8730
rect 1104 8656 15088 8678
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7466 8616 7472 8628
rect 6972 8588 7472 8616
rect 6972 8576 6978 8588
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 11238 8616 11244 8628
rect 10704 8588 11244 8616
rect 10704 8489 10732 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 11716 8548 11744 8579
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13228 8588 13461 8616
rect 13228 8576 13234 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 10888 8520 11744 8548
rect 12253 8551 12311 8557
rect 10888 8489 10916 8520
rect 12253 8517 12265 8551
rect 12299 8548 12311 8551
rect 12434 8548 12440 8560
rect 12299 8520 12440 8548
rect 12299 8517 12311 8520
rect 12253 8511 12311 8517
rect 12434 8508 12440 8520
rect 12492 8548 12498 8560
rect 13538 8548 13544 8560
rect 12492 8520 13544 8548
rect 12492 8508 12498 8520
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14001 8551 14059 8557
rect 14001 8548 14013 8551
rect 13964 8520 14013 8548
rect 13964 8508 13970 8520
rect 14001 8517 14013 8520
rect 14047 8517 14059 8551
rect 14001 8511 14059 8517
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 10612 8412 10640 8443
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 13722 8440 13728 8492
rect 13780 8440 13786 8492
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 10612 8384 11621 8412
rect 10980 8356 11008 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 13587 8415 13645 8421
rect 13587 8412 13599 8415
rect 12400 8384 13599 8412
rect 12400 8372 12406 8384
rect 13587 8381 13599 8384
rect 13633 8381 13645 8415
rect 13587 8375 13645 8381
rect 14090 8372 14096 8424
rect 14148 8372 14154 8424
rect 10962 8304 10968 8356
rect 11020 8304 11026 8356
rect 1104 8186 15088 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 15088 8186
rect 1104 8112 15088 8134
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7432 8044 7849 8072
rect 7432 8032 7438 8044
rect 7837 8041 7849 8044
rect 7883 8072 7895 8075
rect 8202 8072 8208 8084
rect 7883 8044 8208 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7708 7840 7757 7868
rect 7708 7828 7714 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 1104 7642 15088 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 15088 7642
rect 1104 7568 15088 7590
rect 8297 7531 8355 7537
rect 8297 7528 8309 7531
rect 7392 7500 8309 7528
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6236 7432 6653 7460
rect 6236 7420 6242 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 7006 7460 7012 7472
rect 6687 7432 7012 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 7006 7420 7012 7432
rect 7064 7460 7070 7472
rect 7392 7460 7420 7500
rect 8297 7497 8309 7500
rect 8343 7497 8355 7531
rect 8297 7491 8355 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 12529 7531 12587 7537
rect 12529 7528 12541 7531
rect 9732 7500 12541 7528
rect 9732 7488 9738 7500
rect 12529 7497 12541 7500
rect 12575 7497 12587 7531
rect 12529 7491 12587 7497
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 7064 7432 7420 7460
rect 7064 7420 7070 7432
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6328 7364 6837 7392
rect 6328 7352 6334 7364
rect 6825 7361 6837 7364
rect 6871 7392 6883 7395
rect 7190 7392 7196 7404
rect 6871 7364 7196 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7392 7401 7420 7432
rect 7484 7432 8125 7460
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7208 7324 7236 7352
rect 7484 7324 7512 7432
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 8113 7423 8171 7429
rect 11241 7463 11299 7469
rect 11241 7429 11253 7463
rect 11287 7460 11299 7463
rect 11287 7432 11836 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 11330 7352 11336 7404
rect 11388 7352 11394 7404
rect 11808 7401 11836 7432
rect 13538 7401 13544 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 13521 7395 13544 7401
rect 13521 7361 13533 7395
rect 13521 7355 13544 7361
rect 13538 7352 13544 7355
rect 13596 7352 13602 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13722 7392 13728 7404
rect 13679 7364 13728 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 7208 7296 7512 7324
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 13906 7284 13912 7336
rect 13964 7284 13970 7336
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14090 7324 14096 7336
rect 14047 7296 14096 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 6972 7228 7021 7256
rect 6972 7216 6978 7228
rect 7009 7225 7021 7228
rect 7055 7256 7067 7259
rect 7558 7256 7564 7268
rect 7055 7228 7564 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 7340 7160 7389 7188
rect 7340 7148 7346 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7708 7160 8309 7188
rect 7708 7148 7714 7160
rect 8297 7157 8309 7160
rect 8343 7188 8355 7191
rect 8386 7188 8392 7200
rect 8343 7160 8392 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 9766 7188 9772 7200
rect 8527 7160 9772 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 13228 7160 13369 7188
rect 13228 7148 13234 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13357 7151 13415 7157
rect 1104 7098 15088 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 15088 7098
rect 1104 7024 15088 7046
rect 6178 6944 6184 6996
rect 6236 6944 6242 6996
rect 8386 6944 8392 6996
rect 8444 6944 8450 6996
rect 9766 6984 9772 6996
rect 9508 6956 9772 6984
rect 6716 6851 6774 6857
rect 6716 6848 6728 6851
rect 6656 6820 6728 6848
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5491 6752 6285 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6656 6780 6684 6820
rect 6716 6817 6728 6820
rect 6762 6848 6774 6851
rect 6822 6848 6828 6860
rect 6762 6820 6828 6848
rect 6762 6817 6774 6820
rect 6716 6811 6774 6817
rect 6822 6808 6828 6820
rect 6880 6848 6886 6860
rect 6880 6820 7420 6848
rect 6880 6808 6886 6820
rect 6273 6743 6331 6749
rect 6380 6752 6684 6780
rect 5184 6712 5212 6743
rect 6380 6712 6408 6752
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7392 6789 7420 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9508 6857 9536 6956
rect 9766 6944 9772 6956
rect 9824 6984 9830 6996
rect 9824 6956 10180 6984
rect 9824 6944 9830 6956
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 8260 6820 9413 6848
rect 8260 6808 8266 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 10152 6848 10180 6956
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 11388 6956 11437 6984
rect 11388 6944 11394 6956
rect 11425 6953 11437 6956
rect 11471 6984 11483 6987
rect 13722 6984 13728 6996
rect 11471 6956 13728 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 10962 6848 10968 6860
rect 10152 6820 10968 6848
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7742 6780 7748 6792
rect 7699 6752 7748 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 5184 6684 6408 6712
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6681 6515 6715
rect 7282 6712 7288 6724
rect 6457 6675 6515 6681
rect 6840 6684 7288 6712
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6472 6644 6500 6675
rect 6840 6653 6868 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 7392 6712 7420 6743
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9600 6780 9628 6808
rect 10152 6789 10180 6820
rect 10962 6808 10968 6820
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6848 11115 6851
rect 11103 6820 11468 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 9355 6752 9628 6780
rect 9677 6783 9735 6789
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 10011 6783 10069 6789
rect 10011 6780 10023 6783
rect 9723 6752 10023 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 9769 6715 9827 6721
rect 9769 6712 9781 6715
rect 7392 6684 9781 6712
rect 9769 6681 9781 6684
rect 9815 6681 9827 6715
rect 9876 6712 9904 6752
rect 10011 6749 10023 6752
rect 10057 6749 10069 6783
rect 10011 6743 10069 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10376 6752 10425 6780
rect 10376 6740 10382 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11146 6780 11152 6792
rect 10919 6752 11152 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11146 6740 11152 6752
rect 11204 6780 11210 6792
rect 11440 6789 11468 6820
rect 12452 6789 12480 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 12618 6857 12624 6860
rect 12575 6851 12624 6857
rect 12575 6817 12587 6851
rect 12621 6817 12624 6851
rect 12575 6811 12624 6817
rect 12618 6808 12624 6811
rect 12676 6808 12682 6860
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 11204 6752 11253 6780
rect 11204 6740 11210 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12437 6743 12495 6749
rect 12544 6752 12909 6780
rect 11054 6712 11060 6724
rect 9876 6684 11060 6712
rect 9769 6675 9827 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 12069 6715 12127 6721
rect 12069 6681 12081 6715
rect 12115 6681 12127 6715
rect 12069 6675 12127 6681
rect 6236 6616 6500 6644
rect 6825 6647 6883 6653
rect 6236 6604 6242 6616
rect 6825 6613 6837 6647
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 9030 6604 9036 6656
rect 9088 6604 9094 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 10502 6644 10508 6656
rect 9272 6616 10508 6644
rect 9272 6604 9278 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 12084 6644 12112 6675
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 12544 6644 12572 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13173 6753 13231 6759
rect 10652 6616 12572 6644
rect 10652 6604 10658 6616
rect 12710 6604 12716 6656
rect 12768 6604 12774 6656
rect 12912 6644 12940 6743
rect 13173 6724 13185 6753
rect 13219 6724 13231 6753
rect 13170 6672 13176 6724
rect 13228 6672 13234 6724
rect 14090 6712 14096 6724
rect 13280 6684 14096 6712
rect 13078 6644 13084 6656
rect 12912 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6644 13142 6656
rect 13280 6644 13308 6684
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 13136 6616 13308 6644
rect 13136 6604 13142 6616
rect 13906 6604 13912 6656
rect 13964 6604 13970 6656
rect 1104 6554 15088 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 15088 6554
rect 1104 6480 15088 6502
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6440 6334 6452
rect 6638 6440 6644 6452
rect 6328 6412 6644 6440
rect 6328 6400 6334 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 6822 6400 6828 6452
rect 6880 6400 6886 6452
rect 7742 6400 7748 6452
rect 7800 6400 7806 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 11514 6440 11520 6452
rect 10643 6412 11520 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 14090 6440 14096 6452
rect 12216 6412 14096 6440
rect 12216 6400 12222 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 6840 6372 6868 6400
rect 7006 6372 7012 6384
rect 5184 6344 6868 6372
rect 6932 6344 7012 6372
rect 5184 6313 5212 6344
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 6733 6307 6791 6313
rect 5491 6276 6408 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 6380 6177 6408 6276
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 6932 6304 6960 6344
rect 7006 6332 7012 6344
rect 7064 6372 7070 6384
rect 11146 6372 11152 6384
rect 7064 6344 11152 6372
rect 7064 6332 7070 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 6779 6276 6960 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 9030 6304 9036 6316
rect 7883 6276 9036 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6696 6208 6929 6236
rect 6696 6196 6702 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 7484 6236 7512 6267
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9732 6276 9781 6304
rect 9732 6264 9738 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10318 6304 10324 6316
rect 9907 6276 10324 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10594 6304 10600 6316
rect 10459 6276 10600 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 12768 6276 13369 6304
rect 12768 6264 12774 6276
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 8202 6236 8208 6248
rect 7484 6208 8208 6236
rect 6917 6199 6975 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 6365 6171 6423 6177
rect 6365 6137 6377 6171
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 14090 6128 14096 6180
rect 14148 6128 14154 6180
rect 1104 6010 15088 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 15088 6010
rect 1104 5936 15088 5958
rect 1104 5466 15088 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 15088 5466
rect 1104 5392 15088 5414
rect 10686 5312 10692 5364
rect 10744 5312 10750 5364
rect 11146 5312 11152 5364
rect 11204 5312 11210 5364
rect 10597 5287 10655 5293
rect 10597 5253 10609 5287
rect 10643 5284 10655 5287
rect 11698 5284 11704 5296
rect 10643 5256 11704 5284
rect 10643 5253 10655 5256
rect 10597 5247 10655 5253
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 11333 5151 11391 5157
rect 11333 5148 11345 5151
rect 9732 5120 11345 5148
rect 9732 5108 9738 5120
rect 11333 5117 11345 5120
rect 11379 5117 11391 5151
rect 11333 5111 11391 5117
rect 1104 4922 15088 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 15088 4922
rect 1104 4848 15088 4870
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11698 4808 11704 4820
rect 11379 4780 11704 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 11517 4743 11575 4749
rect 11517 4740 11529 4743
rect 11112 4712 11529 4740
rect 11112 4700 11118 4712
rect 11517 4709 11529 4712
rect 11563 4709 11575 4743
rect 11517 4703 11575 4709
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10778 4672 10784 4684
rect 9732 4644 9812 4672
rect 9732 4632 9738 4644
rect 9784 4613 9812 4644
rect 10060 4644 10784 4672
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 9674 4496 9680 4548
rect 9732 4496 9738 4548
rect 9784 4536 9812 4567
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10060 4613 10088 4644
rect 10778 4632 10784 4644
rect 10836 4672 10842 4684
rect 10873 4675 10931 4681
rect 10873 4672 10885 4675
rect 10836 4644 10885 4672
rect 10836 4632 10842 4644
rect 10873 4641 10885 4644
rect 10919 4641 10931 4675
rect 12802 4672 12808 4684
rect 10873 4635 10931 4641
rect 10980 4644 12808 4672
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9916 4576 10057 4604
rect 9916 4564 9922 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 10980 4613 11008 4644
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 10744 4576 10977 4604
rect 10744 4564 10750 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 9950 4536 9956 4548
rect 9784 4508 9956 4536
rect 9950 4496 9956 4508
rect 10008 4536 10014 4548
rect 11348 4536 11376 4567
rect 10008 4508 11376 4536
rect 10008 4496 10014 4508
rect 1104 4378 15088 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 15088 4378
rect 1104 4304 15088 4326
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9208 4267 9266 4273
rect 9208 4264 9220 4267
rect 8996 4236 9220 4264
rect 8996 4224 9002 4236
rect 9208 4233 9220 4236
rect 9254 4264 9266 4267
rect 10226 4264 10232 4276
rect 9254 4236 10232 4264
rect 9254 4233 9266 4236
rect 9208 4227 9266 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 10244 4196 10272 4224
rect 10244 4168 10824 4196
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9214 4128 9220 4140
rect 8895 4100 9220 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 8680 4060 8708 4091
rect 9214 4088 9220 4100
rect 9272 4128 9278 4140
rect 9585 4131 9643 4137
rect 9272 4100 9444 4128
rect 9272 4088 9278 4100
rect 8754 4060 8760 4072
rect 8680 4032 8760 4060
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 9416 4060 9444 4100
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 9766 4128 9772 4140
rect 9631 4100 9772 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10226 4088 10232 4140
rect 10284 4088 10290 4140
rect 10796 4137 10824 4168
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10459 4100 10701 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 10827 4100 13553 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 8812 4032 9260 4060
rect 9416 4032 10088 4060
rect 8812 4020 8818 4032
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 8846 3992 8852 4004
rect 8619 3964 8852 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9232 3992 9260 4032
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 9232 3964 9781 3992
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 9122 3924 9128 3936
rect 9079 3896 9128 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9232 3933 9260 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 10060 3992 10088 4032
rect 10134 4020 10140 4072
rect 10192 4020 10198 4072
rect 10428 3992 10456 4091
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 13188 4001 13216 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 13814 4088 13820 4140
rect 13872 4088 13878 4140
rect 13446 4020 13452 4072
rect 13504 4020 13510 4072
rect 10060 3964 10456 3992
rect 13173 3995 13231 4001
rect 9769 3955 9827 3961
rect 13173 3961 13185 3995
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 9217 3927 9275 3933
rect 9217 3893 9229 3927
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 13262 3884 13268 3936
rect 13320 3884 13326 3936
rect 1104 3834 15088 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 15088 3834
rect 1104 3760 15088 3782
rect 8665 3723 8723 3729
rect 8665 3689 8677 3723
rect 8711 3720 8723 3723
rect 10226 3720 10232 3732
rect 8711 3692 10232 3720
rect 8711 3689 8723 3692
rect 8665 3683 8723 3689
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 8588 3380 8616 3479
rect 8754 3476 8760 3528
rect 8812 3476 8818 3528
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 9140 3525 9168 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10778 3720 10784 3732
rect 10735 3692 10784 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 13814 3720 13820 3732
rect 11756 3692 13820 3720
rect 11756 3680 11762 3692
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14182 3680 14188 3732
rect 14240 3680 14246 3732
rect 9674 3612 9680 3664
rect 9732 3612 9738 3664
rect 9692 3584 9720 3612
rect 9232 3556 9720 3584
rect 12253 3587 12311 3593
rect 9232 3525 9260 3556
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 12299 3556 12449 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12437 3553 12449 3556
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9326 3519 9384 3525
rect 9326 3485 9338 3519
rect 9372 3516 9384 3519
rect 9585 3519 9643 3525
rect 9372 3488 9444 3516
rect 9372 3485 9384 3488
rect 9326 3479 9384 3485
rect 9416 3380 9444 3488
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9631 3488 9689 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10134 3516 10140 3528
rect 9999 3488 10140 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 12342 3476 12348 3528
rect 12400 3476 12406 3528
rect 12704 3519 12762 3525
rect 12704 3485 12716 3519
rect 12750 3516 12762 3519
rect 13446 3516 13452 3528
rect 12750 3488 13452 3516
rect 12750 3485 12762 3488
rect 12704 3479 12762 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13780 3488 14289 3516
rect 13780 3476 13786 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 9858 3380 9864 3392
rect 8588 3352 9864 3380
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 1104 3290 15088 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 15088 3290
rect 1104 3216 15088 3238
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 12860 3148 14381 3176
rect 12860 3136 12866 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 14369 3139 14427 3145
rect 13262 3117 13268 3120
rect 13256 3108 13268 3117
rect 13223 3080 13268 3108
rect 13256 3071 13268 3080
rect 13262 3068 13268 3071
rect 13320 3068 13326 3120
rect 8846 3000 8852 3052
rect 8904 3000 8910 3052
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12400 2944 13001 2972
rect 12400 2932 12406 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 9858 2796 9864 2848
rect 9916 2796 9922 2848
rect 1104 2746 15088 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 15088 2746
rect 1104 2672 15088 2694
rect 1104 2202 15088 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 15088 2202
rect 1104 2128 15088 2150
<< via1 >>
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 14004 15079 14056 15088
rect 14004 15045 14013 15079
rect 14013 15045 14047 15079
rect 14047 15045 14056 15079
rect 14004 15036 14056 15045
rect 13728 15011 13780 15020
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 12164 14900 12216 14952
rect 13084 14832 13136 14884
rect 13176 14764 13228 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 9312 14560 9364 14612
rect 12164 14560 12216 14612
rect 14004 14560 14056 14612
rect 10692 14535 10744 14544
rect 10692 14501 10701 14535
rect 10701 14501 10735 14535
rect 10735 14501 10744 14535
rect 10692 14492 10744 14501
rect 11060 14492 11112 14544
rect 4620 14356 4672 14408
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 13084 14356 13136 14408
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 9772 14288 9824 14340
rect 10876 14288 10928 14340
rect 7564 14220 7616 14272
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 5448 13948 5500 14000
rect 12624 14016 12676 14068
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 4620 13812 4672 13864
rect 6736 13855 6788 13864
rect 6736 13821 6745 13855
rect 6745 13821 6779 13855
rect 6779 13821 6788 13855
rect 6736 13812 6788 13821
rect 6460 13744 6512 13796
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9220 13948 9272 14000
rect 9312 13991 9364 14000
rect 9312 13957 9321 13991
rect 9321 13957 9355 13991
rect 9355 13957 9364 13991
rect 9312 13948 9364 13957
rect 13452 13948 13504 14000
rect 7656 13880 7708 13932
rect 8668 13880 8720 13932
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 7840 13812 7892 13864
rect 7932 13855 7984 13864
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 8484 13812 8536 13864
rect 6920 13676 6972 13728
rect 8392 13744 8444 13796
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 7472 13676 7524 13728
rect 10508 13880 10560 13932
rect 12440 13880 12492 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 10232 13676 10284 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 6828 13472 6880 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13360 13472 13412 13524
rect 6460 13447 6512 13456
rect 6460 13413 6469 13447
rect 6469 13413 6503 13447
rect 6503 13413 6512 13447
rect 6460 13404 6512 13413
rect 6920 13404 6972 13456
rect 7012 13404 7064 13456
rect 7288 13336 7340 13388
rect 8024 13336 8076 13388
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 6552 13268 6604 13320
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 7840 13268 7892 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 8484 13268 8536 13320
rect 10876 13336 10928 13388
rect 11704 13336 11756 13388
rect 12624 13379 12676 13388
rect 12624 13345 12647 13379
rect 12647 13345 12676 13379
rect 12624 13336 12676 13345
rect 6552 13132 6604 13184
rect 6644 13132 6696 13184
rect 7472 13200 7524 13252
rect 7932 13132 7984 13184
rect 10232 13268 10284 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 14096 13336 14148 13388
rect 11152 13200 11204 13252
rect 11428 13200 11480 13252
rect 12256 13200 12308 13252
rect 13728 13268 13780 13320
rect 12992 13243 13044 13252
rect 12992 13209 13001 13243
rect 13001 13209 13035 13243
rect 13035 13209 13044 13243
rect 12992 13200 13044 13209
rect 13084 13243 13136 13252
rect 13084 13209 13093 13243
rect 13093 13209 13127 13243
rect 13127 13209 13136 13243
rect 13084 13200 13136 13209
rect 11244 13175 11296 13184
rect 11244 13141 11253 13175
rect 11253 13141 11287 13175
rect 11287 13141 11296 13175
rect 11244 13132 11296 13141
rect 12716 13132 12768 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 6552 12928 6604 12980
rect 8024 12928 8076 12980
rect 5908 12860 5960 12912
rect 7012 12903 7064 12912
rect 7012 12869 7021 12903
rect 7021 12869 7055 12903
rect 7055 12869 7064 12903
rect 7012 12860 7064 12869
rect 7840 12860 7892 12912
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 7380 12792 7432 12844
rect 7564 12792 7616 12844
rect 11428 12792 11480 12844
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 6828 12724 6880 12776
rect 8484 12656 8536 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 6828 12384 6880 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 13452 12427 13504 12436
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 14188 12248 14240 12300
rect 6920 12180 6972 12232
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 10324 12180 10376 12232
rect 13912 12223 13964 12232
rect 13912 12189 13921 12223
rect 13921 12189 13955 12223
rect 13955 12189 13964 12223
rect 13912 12180 13964 12189
rect 13820 12112 13872 12164
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 7472 11092 7524 11144
rect 9772 11092 9824 11144
rect 10140 11092 10192 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 12716 11092 12768 11144
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 5908 10956 5960 11008
rect 6736 11024 6788 11076
rect 10968 10999 11020 11008
rect 10968 10965 10977 10999
rect 10977 10965 11011 10999
rect 11011 10965 11020 10999
rect 10968 10956 11020 10965
rect 12348 10956 12400 11008
rect 13544 10999 13596 11008
rect 13544 10965 13553 10999
rect 13553 10965 13587 10999
rect 13587 10965 13596 10999
rect 13544 10956 13596 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5908 10795 5960 10804
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 4620 10616 4672 10668
rect 5724 10616 5776 10668
rect 6092 10412 6144 10464
rect 7012 10752 7064 10804
rect 8024 10752 8076 10804
rect 10968 10752 11020 10804
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7932 10684 7984 10736
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 10232 10684 10284 10736
rect 11244 10684 11296 10736
rect 6828 10548 6880 10600
rect 7380 10548 7432 10600
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 7656 10412 7708 10464
rect 9864 10548 9916 10600
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 10876 10616 10928 10668
rect 13728 10684 13780 10736
rect 14556 10727 14608 10736
rect 14556 10693 14565 10727
rect 14565 10693 14599 10727
rect 14599 10693 14608 10727
rect 14556 10684 14608 10693
rect 12716 10548 12768 10600
rect 9496 10412 9548 10464
rect 14372 10548 14424 10600
rect 14556 10480 14608 10532
rect 14096 10412 14148 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 6276 10208 6328 10260
rect 7656 10208 7708 10260
rect 8024 10208 8076 10260
rect 12808 10208 12860 10260
rect 4620 10140 4672 10192
rect 8392 10140 8444 10192
rect 10876 10140 10928 10192
rect 6092 10072 6144 10124
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7380 10072 7432 10124
rect 7104 9979 7156 9988
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 7196 9868 7248 9920
rect 7840 10004 7892 10056
rect 8116 10072 8168 10124
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 10232 10072 10284 10124
rect 13544 10072 13596 10124
rect 7564 9936 7616 9988
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 10968 10004 11020 10056
rect 13084 10047 13136 10056
rect 13084 10013 13107 10047
rect 13107 10013 13136 10047
rect 13084 10004 13136 10013
rect 13728 10004 13780 10056
rect 12716 9936 12768 9988
rect 14096 9936 14148 9988
rect 7932 9868 7984 9920
rect 11244 9868 11296 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 6000 9664 6052 9716
rect 6552 9639 6604 9648
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 7932 9664 7984 9716
rect 7472 9596 7524 9648
rect 9680 9596 9732 9648
rect 10968 9596 11020 9648
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 6828 9503 6880 9512
rect 6828 9469 6854 9503
rect 6854 9469 6880 9503
rect 6828 9460 6880 9469
rect 4712 9324 4764 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 4620 8916 4672 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 7380 9052 7432 9104
rect 6920 8984 6972 9036
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 7564 8916 7616 8968
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 6920 8891 6972 8900
rect 6920 8857 6929 8891
rect 6929 8857 6963 8891
rect 6963 8857 6972 8891
rect 6920 8848 6972 8857
rect 12624 8848 12676 8900
rect 13176 8959 13228 8968
rect 13176 8925 13185 8959
rect 13185 8925 13219 8959
rect 13219 8925 13228 8959
rect 13176 8916 13228 8925
rect 14096 8848 14148 8900
rect 12440 8780 12492 8832
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 6920 8576 6972 8628
rect 7472 8576 7524 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 11244 8576 11296 8628
rect 13176 8576 13228 8628
rect 12440 8508 12492 8560
rect 13544 8508 13596 8560
rect 13912 8508 13964 8560
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 12348 8372 12400 8424
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 10968 8304 11020 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 7380 8032 7432 8084
rect 8208 8032 8260 8084
rect 7656 7828 7708 7880
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 6184 7420 6236 7472
rect 7012 7420 7064 7472
rect 9680 7488 9732 7540
rect 6276 7352 6328 7404
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 13544 7395 13596 7404
rect 13544 7361 13567 7395
rect 13567 7361 13596 7395
rect 13544 7352 13596 7361
rect 13728 7352 13780 7404
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 14096 7284 14148 7336
rect 6920 7216 6972 7268
rect 7564 7216 7616 7268
rect 7288 7148 7340 7200
rect 7656 7148 7708 7200
rect 8392 7148 8444 7200
rect 9772 7148 9824 7200
rect 13176 7148 13228 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 6828 6808 6880 6860
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 8208 6808 8260 6860
rect 9772 6944 9824 6996
rect 9588 6808 9640 6860
rect 11336 6944 11388 6996
rect 6184 6604 6236 6656
rect 7288 6672 7340 6724
rect 7748 6740 7800 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 10968 6808 11020 6860
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10324 6740 10376 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11152 6740 11204 6792
rect 13728 6944 13780 6996
rect 12624 6808 12676 6860
rect 11060 6672 11112 6724
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 9220 6604 9272 6656
rect 10508 6604 10560 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 10600 6604 10652 6613
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 13176 6719 13185 6724
rect 13185 6719 13219 6724
rect 13219 6719 13228 6724
rect 13176 6672 13228 6719
rect 13084 6604 13136 6656
rect 14096 6672 14148 6724
rect 13912 6647 13964 6656
rect 13912 6613 13921 6647
rect 13921 6613 13955 6647
rect 13955 6613 13964 6647
rect 13912 6604 13964 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 6276 6400 6328 6452
rect 6644 6400 6696 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7748 6443 7800 6452
rect 7748 6409 7757 6443
rect 7757 6409 7791 6443
rect 7791 6409 7800 6443
rect 7748 6400 7800 6409
rect 11520 6400 11572 6452
rect 12164 6400 12216 6452
rect 14096 6400 14148 6452
rect 7012 6332 7064 6384
rect 11152 6332 11204 6384
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 6644 6196 6696 6248
rect 9036 6264 9088 6316
rect 9680 6264 9732 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10600 6264 10652 6316
rect 12716 6264 12768 6316
rect 8208 6196 8260 6248
rect 13084 6239 13136 6248
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 14096 6171 14148 6180
rect 14096 6137 14105 6171
rect 14105 6137 14139 6171
rect 14139 6137 14148 6171
rect 14096 6128 14148 6137
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 11704 5244 11756 5296
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 9680 5108 9732 5160
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 11704 4768 11756 4820
rect 11060 4700 11112 4752
rect 9680 4632 9732 4684
rect 9680 4539 9732 4548
rect 9680 4505 9689 4539
rect 9689 4505 9723 4539
rect 9723 4505 9732 4539
rect 9680 4496 9732 4505
rect 9864 4564 9916 4616
rect 10784 4632 10836 4684
rect 10692 4564 10744 4616
rect 12808 4632 12860 4684
rect 9956 4496 10008 4548
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 8944 4224 8996 4276
rect 10232 4224 10284 4276
rect 9220 4088 9272 4140
rect 8760 4020 8812 4072
rect 9772 4088 9824 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 8852 3952 8904 4004
rect 9128 3884 9180 3936
rect 10140 4063 10192 4072
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 10140 4020 10192 4029
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 10232 3680 10284 3732
rect 10784 3680 10836 3732
rect 11704 3680 11756 3732
rect 13820 3723 13872 3732
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 9680 3612 9732 3664
rect 10140 3476 10192 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 13452 3476 13504 3528
rect 13728 3476 13780 3528
rect 9864 3340 9916 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 12808 3136 12860 3188
rect 13268 3111 13320 3120
rect 13268 3077 13302 3111
rect 13302 3077 13320 3111
rect 13268 3068 13320 3077
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 12348 2932 12400 2984
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 11058 16416 11114 16425
rect 11058 16351 11114 16360
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 4632 13870 4660 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 10674 4660 13806
rect 5460 13530 5488 13942
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5920 12918 5948 14350
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7380 13932 7432 13938
rect 7432 13892 7512 13920
rect 7380 13874 7432 13880
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6472 13462 6500 13738
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 13190 6592 13262
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6564 12986 6592 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 6656 12850 6684 13126
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6748 12782 6776 13806
rect 6932 13734 6960 13806
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 12782 6868 13466
rect 6932 13462 6960 13670
rect 7024 13462 7052 13806
rect 7484 13734 7512 13892
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12442 6868 12718
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5920 10810 5948 10950
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6748 10674 6776 11018
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10198 4660 10610
rect 5736 10266 5764 10610
rect 6840 10606 6868 12378
rect 6932 12238 6960 13398
rect 7024 12918 7052 13398
rect 7300 13394 7328 13670
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7484 13258 7512 13670
rect 7576 13326 7604 14214
rect 9232 14006 9260 14350
rect 9324 14006 9352 14554
rect 11072 14550 11100 16351
rect 14002 15736 14058 15745
rect 14002 15671 14058 15680
rect 14016 15094 14044 15671
rect 14004 15088 14056 15094
rect 13910 15056 13966 15065
rect 13728 15020 13780 15026
rect 14004 15030 14056 15036
rect 13910 14991 13966 15000
rect 13728 14962 13780 14968
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12176 14618 12204 14894
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 10674 6960 12174
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8974 4660 10134
rect 6104 10130 6132 10406
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6288 10062 6316 10202
rect 6840 10130 6868 10542
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 6012 9722 6040 9998
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6932 9874 6960 10610
rect 7024 10062 7052 10746
rect 7392 10606 7420 12786
rect 7484 11150 7512 13194
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 10130 7420 10542
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6564 9654 6592 9862
rect 6932 9846 7052 9874
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8974 4752 9318
rect 6840 9178 6868 9454
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 9042 6960 9658
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 6932 8634 6960 8842
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 7024 7478 7052 9846
rect 7116 9586 7144 9930
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 6196 7002 6224 7414
rect 7208 7410 7236 9862
rect 7392 9110 7420 10066
rect 7484 9654 7512 11086
rect 7668 10674 7696 13874
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 7852 13326 7880 13806
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7852 12918 7880 13262
rect 7944 13190 7972 13806
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7852 12238 7880 12854
rect 7944 12442 7972 13126
rect 8036 12986 8064 13330
rect 8404 13326 8432 13738
rect 8496 13326 8524 13806
rect 8680 13530 8708 13874
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 9784 13394 9812 14282
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13938 10548 14214
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7668 10470 7696 10610
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10266 7696 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7392 8090 7420 9046
rect 7484 8634 7512 9590
rect 7576 8974 7604 9930
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6196 6662 6224 6938
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 6288 6458 6316 7346
rect 7576 7274 7604 8910
rect 7668 7886 7696 10202
rect 7852 10062 7880 12174
rect 7944 10742 7972 12378
rect 8036 10826 8064 12922
rect 8496 12714 8524 13262
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 9784 11150 9812 13330
rect 10244 13326 10272 13670
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 8036 10810 8156 10826
rect 8024 10804 8156 10810
rect 8076 10798 8156 10804
rect 8024 10746 8076 10752
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7944 9926 7972 10542
rect 8036 10266 8064 10610
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8128 10130 8156 10798
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 8404 10198 8432 10542
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 9508 10130 9536 10406
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9876 10062 9904 10542
rect 10060 10062 10088 10542
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 9722 7972 9862
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 9692 9654 9720 9998
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6458 6868 6802
rect 6932 6798 6960 7210
rect 7668 7206 7696 7822
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6656 6254 6684 6394
rect 7024 6390 7052 6734
rect 7300 6730 7328 7142
rect 8220 6866 8248 8026
rect 9692 7546 9720 9590
rect 10152 9042 10180 11086
rect 10244 10742 10272 11086
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10244 10130 10272 10542
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 7002 8432 7142
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 9588 6860 9640 6866
rect 9692 6848 9720 7482
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 7002 9812 7142
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 10336 6882 10364 12174
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8634 10456 8910
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 9640 6820 9720 6848
rect 9588 6802 9640 6808
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7300 6322 7328 6666
rect 7760 6458 7788 6734
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 8220 6254 8248 6802
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6662 9260 6734
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9048 6322 9076 6598
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8772 3534 8800 4014
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 8864 3058 8892 3946
rect 8956 3534 8984 4218
rect 9232 4146 9260 6598
rect 9692 6322 9720 6820
rect 10244 6854 10364 6882
rect 10244 6798 10272 6854
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9692 5166 9720 6258
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 4690 9720 5102
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9140 3058 9168 3878
rect 9692 3670 9720 4490
rect 9876 4146 9904 4558
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9968 4146 9996 4490
rect 10244 4282 10272 6734
rect 10336 6322 10364 6734
rect 10520 6662 10548 6734
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6322 10640 6598
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10704 5370 10732 14486
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10888 13394 10916 14282
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 11256 13326 11284 13670
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11164 12434 11192 13194
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11072 12406 11192 12434
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 10810 11008 10950
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10198 10916 10610
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10980 10062 11008 10746
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 8498 11008 9590
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 6866 11008 8298
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11072 6730 11100 12406
rect 11256 10742 11284 13126
rect 11440 12850 11468 13194
rect 11716 13025 11744 13330
rect 11702 13016 11758 13025
rect 11702 12951 11758 12960
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 9926 11284 10678
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 8634 11284 9862
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11716 8498 11744 12951
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11348 7002 11376 7346
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10704 4622 10732 5306
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10796 4690 10824 5170
rect 11072 4758 11100 6666
rect 11164 6390 11192 6734
rect 11532 6458 11560 7278
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11164 5370 11192 6326
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11716 5302 11744 8434
rect 12176 7426 12204 14554
rect 13096 14414 13124 14826
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14414 13216 14758
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12452 13530 12480 13874
rect 12636 13705 12664 14010
rect 13096 13870 13124 14350
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12992 13728 13044 13734
rect 12622 13696 12678 13705
rect 12992 13670 13044 13676
rect 12622 13631 12678 13640
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12636 13394 12664 13631
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 13004 13258 13032 13670
rect 13096 13258 13124 13806
rect 13372 13530 13400 13874
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12268 7585 12296 13194
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 11150 12756 13126
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 8430 12388 10950
rect 12728 10606 12756 11086
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 9994 12756 10542
rect 12820 10266 12848 11086
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8566 12480 8774
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12254 7576 12310 7585
rect 12254 7511 12310 7520
rect 12176 7398 12296 7426
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6458 12204 6666
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11716 4826 11744 5238
rect 12268 4865 12296 7398
rect 12360 5545 12388 8366
rect 12636 6905 12664 8842
rect 12622 6896 12678 6905
rect 12622 6831 12624 6840
rect 12676 6831 12678 6840
rect 12624 6802 12676 6808
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6322 12756 6598
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12346 5536 12402 5545
rect 12346 5471 12402 5480
rect 12254 4856 12310 4865
rect 11704 4820 11756 4826
rect 12254 4791 12310 4800
rect 11704 4762 11756 4768
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9784 4026 9812 4082
rect 10140 4072 10192 4078
rect 9784 3998 9904 4026
rect 10140 4014 10192 4020
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9876 3398 9904 3998
rect 10152 3534 10180 4014
rect 10244 3738 10272 4082
rect 10796 3738 10824 4626
rect 11716 3738 11744 4762
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12820 4078 12848 4626
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9876 2854 9904 3334
rect 12360 2990 12388 3470
rect 12820 3194 12848 4014
rect 13004 3505 13032 13194
rect 13464 12442 13492 13942
rect 13740 13326 13768 14962
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13544 11008 13596 11014
rect 13542 10976 13544 10985
rect 13596 10976 13598 10985
rect 13542 10911 13598 10920
rect 13556 10130 13584 10911
rect 13740 10742 13768 13262
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 13832 12170 13860 12271
rect 13924 12238 13952 14991
rect 14016 14618 14044 15030
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14094 14376 14150 14385
rect 14094 14311 14150 14320
rect 14108 14074 14136 14311
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14108 13394 14136 14010
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13740 10062 13768 10678
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13096 9625 13124 9998
rect 13082 9616 13138 9625
rect 13082 9551 13138 9560
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8634 13216 8910
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13556 8265 13584 8502
rect 13740 8498 13768 9998
rect 14108 9994 14136 10406
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13910 8936 13966 8945
rect 14108 8906 14136 9930
rect 13910 8871 13966 8880
rect 14096 8900 14148 8906
rect 13924 8838 13952 8871
rect 14096 8842 14148 8848
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8566 13952 8774
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13542 8256 13598 8265
rect 13542 8191 13598 8200
rect 13556 7410 13584 8191
rect 13740 7410 13768 8434
rect 14108 8430 14136 8842
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6730 13216 7142
rect 13740 7002 13768 7346
rect 14108 7342 14136 8366
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13924 6662 13952 7278
rect 14108 6730 14136 7278
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13096 6254 13124 6598
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13924 4185 13952 6598
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14108 6225 14136 6394
rect 14094 6216 14150 6225
rect 14094 6151 14096 6160
rect 14148 6151 14150 6160
rect 14096 6122 14148 6128
rect 13910 4176 13966 4185
rect 13820 4140 13872 4146
rect 13910 4111 13966 4120
rect 13820 4082 13872 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12990 3496 13046 3505
rect 12990 3431 13046 3440
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13280 3126 13308 3878
rect 13464 3534 13492 4014
rect 13832 3738 13860 4082
rect 14200 3738 14228 12242
rect 14554 11656 14610 11665
rect 14554 11591 14610 11600
rect 14568 10742 14596 11591
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10305 14412 10542
rect 14568 10538 14596 10678
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14370 10296 14426 10305
rect 14370 10231 14426 10240
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 9864 2848 9916 2854
rect 9862 2816 9864 2825
rect 9916 2816 9918 2825
rect 4214 2748 4522 2757
rect 9862 2751 9918 2760
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 12360 1465 12388 2926
rect 13740 2145 13768 3470
rect 13726 2136 13782 2145
rect 13726 2071 13782 2080
rect 12346 1456 12402 1465
rect 12346 1391 12402 1400
<< via2 >>
rect 11058 16360 11114 16416
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 14002 15680 14058 15736
rect 13910 15000 13966 15056
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 11702 12960 11758 13016
rect 12622 13640 12678 13696
rect 12254 7520 12310 7576
rect 12622 6860 12678 6896
rect 12622 6840 12624 6860
rect 12624 6840 12676 6860
rect 12676 6840 12678 6860
rect 12346 5480 12402 5536
rect 12254 4800 12310 4856
rect 13542 10956 13544 10976
rect 13544 10956 13596 10976
rect 13596 10956 13598 10976
rect 13542 10920 13598 10956
rect 13818 12280 13874 12336
rect 14094 14320 14150 14376
rect 13082 9560 13138 9616
rect 13910 8880 13966 8936
rect 13542 8200 13598 8256
rect 14094 6180 14150 6216
rect 14094 6160 14096 6180
rect 14096 6160 14148 6180
rect 14148 6160 14150 6180
rect 13910 4120 13966 4176
rect 12990 3440 13046 3496
rect 14554 11600 14610 11656
rect 14370 10240 14426 10296
rect 9862 2796 9864 2816
rect 9864 2796 9916 2816
rect 9916 2796 9918 2816
rect 9862 2760 9918 2796
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 13726 2080 13782 2136
rect 12346 1400 12402 1456
<< metal3 >>
rect 11053 16418 11119 16421
rect 15424 16418 16224 16448
rect 11053 16416 16224 16418
rect 11053 16360 11058 16416
rect 11114 16360 16224 16416
rect 11053 16358 16224 16360
rect 11053 16355 11119 16358
rect 15424 16328 16224 16358
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 13997 15738 14063 15741
rect 15424 15738 16224 15768
rect 13997 15736 16224 15738
rect 13997 15680 14002 15736
rect 14058 15680 16224 15736
rect 13997 15678 16224 15680
rect 13997 15675 14063 15678
rect 15424 15648 16224 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 13905 15058 13971 15061
rect 15424 15058 16224 15088
rect 13905 15056 16224 15058
rect 13905 15000 13910 15056
rect 13966 15000 16224 15056
rect 13905 14998 16224 15000
rect 13905 14995 13971 14998
rect 15424 14968 16224 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 14089 14378 14155 14381
rect 15424 14378 16224 14408
rect 14089 14376 16224 14378
rect 14089 14320 14094 14376
rect 14150 14320 16224 14376
rect 14089 14318 16224 14320
rect 14089 14315 14155 14318
rect 15424 14288 16224 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 12617 13698 12683 13701
rect 15424 13698 16224 13728
rect 12617 13696 16224 13698
rect 12617 13640 12622 13696
rect 12678 13640 16224 13696
rect 12617 13638 16224 13640
rect 12617 13635 12683 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 15424 13608 16224 13638
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 11697 13018 11763 13021
rect 15424 13018 16224 13048
rect 11697 13016 16224 13018
rect 11697 12960 11702 13016
rect 11758 12960 16224 13016
rect 11697 12958 16224 12960
rect 11697 12955 11763 12958
rect 15424 12928 16224 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 13813 12338 13879 12341
rect 15424 12338 16224 12368
rect 13813 12336 16224 12338
rect 13813 12280 13818 12336
rect 13874 12280 16224 12336
rect 13813 12278 16224 12280
rect 13813 12275 13879 12278
rect 15424 12248 16224 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 14549 11658 14615 11661
rect 15424 11658 16224 11688
rect 14549 11656 16224 11658
rect 14549 11600 14554 11656
rect 14610 11600 16224 11656
rect 14549 11598 16224 11600
rect 14549 11595 14615 11598
rect 15424 11568 16224 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 13537 10978 13603 10981
rect 15424 10978 16224 11008
rect 13537 10976 16224 10978
rect 13537 10920 13542 10976
rect 13598 10920 16224 10976
rect 13537 10918 16224 10920
rect 13537 10915 13603 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 15424 10888 16224 10918
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 14365 10298 14431 10301
rect 15424 10298 16224 10328
rect 14365 10296 16224 10298
rect 14365 10240 14370 10296
rect 14426 10240 16224 10296
rect 14365 10238 16224 10240
rect 14365 10235 14431 10238
rect 15424 10208 16224 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 13077 9618 13143 9621
rect 15424 9618 16224 9648
rect 13077 9616 16224 9618
rect 13077 9560 13082 9616
rect 13138 9560 16224 9616
rect 13077 9558 16224 9560
rect 13077 9555 13143 9558
rect 15424 9528 16224 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 13905 8938 13971 8941
rect 15424 8938 16224 8968
rect 13905 8936 16224 8938
rect 13905 8880 13910 8936
rect 13966 8880 16224 8936
rect 13905 8878 16224 8880
rect 13905 8875 13971 8878
rect 15424 8848 16224 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 13537 8258 13603 8261
rect 15424 8258 16224 8288
rect 13537 8256 16224 8258
rect 13537 8200 13542 8256
rect 13598 8200 16224 8256
rect 13537 8198 16224 8200
rect 13537 8195 13603 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 15424 8168 16224 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 12249 7578 12315 7581
rect 15424 7578 16224 7608
rect 12249 7576 16224 7578
rect 12249 7520 12254 7576
rect 12310 7520 16224 7576
rect 12249 7518 16224 7520
rect 12249 7515 12315 7518
rect 15424 7488 16224 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12617 6898 12683 6901
rect 15424 6898 16224 6928
rect 12617 6896 16224 6898
rect 12617 6840 12622 6896
rect 12678 6840 16224 6896
rect 12617 6838 16224 6840
rect 12617 6835 12683 6838
rect 15424 6808 16224 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 14089 6218 14155 6221
rect 15424 6218 16224 6248
rect 14089 6216 16224 6218
rect 14089 6160 14094 6216
rect 14150 6160 16224 6216
rect 14089 6158 16224 6160
rect 14089 6155 14155 6158
rect 15424 6128 16224 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12341 5538 12407 5541
rect 15424 5538 16224 5568
rect 12341 5536 16224 5538
rect 12341 5480 12346 5536
rect 12402 5480 16224 5536
rect 12341 5478 16224 5480
rect 12341 5475 12407 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 15424 5448 16224 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12249 4858 12315 4861
rect 15424 4858 16224 4888
rect 12249 4856 16224 4858
rect 12249 4800 12254 4856
rect 12310 4800 16224 4856
rect 12249 4798 16224 4800
rect 12249 4795 12315 4798
rect 15424 4768 16224 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 13905 4178 13971 4181
rect 15424 4178 16224 4208
rect 13905 4176 16224 4178
rect 13905 4120 13910 4176
rect 13966 4120 16224 4176
rect 13905 4118 16224 4120
rect 13905 4115 13971 4118
rect 15424 4088 16224 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12985 3498 13051 3501
rect 15424 3498 16224 3528
rect 12985 3496 16224 3498
rect 12985 3440 12990 3496
rect 13046 3440 16224 3496
rect 12985 3438 16224 3440
rect 12985 3435 13051 3438
rect 15424 3408 16224 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 9857 2818 9923 2821
rect 15424 2818 16224 2848
rect 9857 2816 16224 2818
rect 9857 2760 9862 2816
rect 9918 2760 16224 2816
rect 9857 2758 16224 2760
rect 9857 2755 9923 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 15424 2728 16224 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 13721 2138 13787 2141
rect 15424 2138 16224 2168
rect 13721 2136 16224 2138
rect 13721 2080 13726 2136
rect 13782 2080 16224 2136
rect 13721 2078 16224 2080
rect 13721 2075 13787 2078
rect 15424 2048 16224 2078
rect 12341 1458 12407 1461
rect 15424 1458 16224 1488
rect 12341 1456 16224 1458
rect 12341 1400 12346 1456
rect 12402 1400 16224 1456
rect 12341 1398 16224 1400
rect 12341 1395 12407 1398
rect 15424 1368 16224 1398
<< via3 >>
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 15808 4528 15824
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 15264 5188 15824
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _067_
timestamp -25199
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp -25199
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp -25199
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp -25199
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp -25199
transform 1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp -25199
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp -25199
transform -1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _074_
timestamp -25199
transform -1 0 13892 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _075_
timestamp -25199
transform -1 0 7636 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _076_
timestamp -25199
transform -1 0 7544 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _077_
timestamp -25199
transform 1 0 6624 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _078_
timestamp -25199
transform 1 0 9752 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _079_
timestamp -25199
transform 1 0 5520 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _080_
timestamp -25199
transform -1 0 11132 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _081_
timestamp -25199
transform 1 0 5336 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_2  _082_
timestamp -25199
transform -1 0 11040 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _083_
timestamp -25199
transform -1 0 11408 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_2  _084_
timestamp -25199
transform 1 0 10764 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _085_
timestamp -25199
transform 1 0 11132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _086_
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _087_
timestamp -25199
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_2  _088_
timestamp -25199
transform -1 0 8372 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _089_
timestamp -25199
transform 1 0 6256 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _090_
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_2  _091_
timestamp -25199
transform 1 0 5612 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _092_
timestamp -25199
transform -1 0 9384 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _093_
timestamp -25199
transform -1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _094_
timestamp -25199
transform -1 0 8832 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_2  _095_
timestamp -25199
transform -1 0 8740 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _096_
timestamp -25199
transform 1 0 8096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _097_
timestamp -25199
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _098_
timestamp -25199
transform -1 0 11592 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp -25199
transform -1 0 11408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _100_
timestamp -25199
transform 1 0 10304 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _101_
timestamp -25199
transform -1 0 10120 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _102_
timestamp -25199
transform -1 0 8924 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _103_
timestamp -25199
transform -1 0 8832 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _104_
timestamp -25199
transform -1 0 10120 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _105_
timestamp -25199
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _106_
timestamp -25199
transform -1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _107_
timestamp -25199
transform -1 0 10580 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _108_
timestamp -25199
transform -1 0 10488 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _109_
timestamp -25199
transform -1 0 11132 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _110_
timestamp -25199
transform 1 0 10212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _111_
timestamp -25199
transform -1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _112_
timestamp -25199
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _113_
timestamp -25199
transform 1 0 13156 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _114_
timestamp -25199
transform -1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _115_
timestamp -25199
transform 1 0 12328 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _116_
timestamp -25199
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _117_
timestamp -25199
transform 1 0 13340 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _118_
timestamp -25199
transform 1 0 13340 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _119_
timestamp -25199
transform 1 0 13248 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _121_
timestamp -25199
transform 1 0 6256 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _122_
timestamp -25199
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _123_
timestamp -25199
transform 1 0 7268 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _124_
timestamp -25199
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _125_
timestamp -25199
transform 1 0 10488 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _126_
timestamp -25199
transform -1 0 7636 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _127_
timestamp -25199
transform -1 0 7176 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_2  _128_
timestamp -25199
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _129_
timestamp -25199
transform -1 0 7176 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _130_
timestamp -25199
transform -1 0 7084 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _131_
timestamp -25199
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _132_
timestamp -25199
transform 1 0 12788 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _133_
timestamp -25199
transform 1 0 13340 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _134_
timestamp -25199
transform 1 0 12420 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _135_
timestamp -25199
transform 1 0 12972 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dlxtn_1  _136_
timestamp -25199
transform 1 0 8832 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _137_
timestamp -25199
transform 1 0 9660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _138_
timestamp -25199
transform 1 0 9844 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dlxtn_1  _139_
timestamp -25199
transform 1 0 9936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _140_
timestamp -25199
transform 1 0 5612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _141_
timestamp -25199
transform 1 0 4416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _142_
timestamp -25199
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _143_
timestamp -25199
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _144_
timestamp -25199
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _145_
timestamp -25199
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _146_
timestamp -25199
transform 1 0 10120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _147_
timestamp -25199
transform 1 0 12512 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _148_
timestamp -25199
transform 1 0 13064 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _149_
timestamp -25199
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _150_
timestamp -25199
transform 1 0 11960 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _151_
timestamp -25199
transform 1 0 12788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _152_
timestamp -25199
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _153_
timestamp -25199
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _154_
timestamp -25199
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _155_
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _156_
timestamp -25199
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _157_
timestamp -25199
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _158_
timestamp -25199
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636943256
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp -25199
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp -25199
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636943256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636943256
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp -25199
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp -25199
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636943256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_81
timestamp -25199
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_96
timestamp 1636943256
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_108
timestamp -25199
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636943256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_125
timestamp -25199
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_146
timestamp -25199
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636943256
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636943256
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636943256
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_77
timestamp -25199
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_105
timestamp 1636943256
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_117
timestamp -25199
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_144
timestamp -25199
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_148
timestamp -25199
transform 1 0 14720 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636943256
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636943256
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp -25199
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp -25199
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_77
timestamp -25199
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp -25199
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636943256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_125
timestamp -25199
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_139
timestamp -25199
transform 1 0 13892 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_147
timestamp -25199
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636943256
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636943256
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636943256
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636943256
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636943256
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp -25199
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp -25199
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_98
timestamp -25199
transform 1 0 10120 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_104
timestamp -25199
transform 1 0 10672 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_115
timestamp 1636943256
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_127
timestamp 1636943256
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp -25199
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp -25199
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636943256
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636943256
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636943256
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636943256
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp -25199
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp -25199
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636943256
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_93
timestamp -25199
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp -25199
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636943256
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636943256
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636943256
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636943256
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636943256
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636943256
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636943256
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636943256
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp -25199
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636943256
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636943256
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636943256
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636943256
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp -25199
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp -25199
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_141
timestamp -25199
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636943256
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636943256
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636943256
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_39
timestamp -25199
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_43
timestamp -25199
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_66
timestamp -25199
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_74
timestamp 1636943256
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_86
timestamp -25199
transform 1 0 9016 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_97
timestamp -25199
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp -25199
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp -25199
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636943256
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_125
timestamp -25199
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_129
timestamp -25199
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_142
timestamp -25199
transform 1 0 14168 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_148
timestamp -25199
transform 1 0 14720 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636943256
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636943256
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp -25199
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636943256
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp -25199
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_65
timestamp -25199
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp -25199
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_114
timestamp -25199
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_118
timestamp -25199
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp -25199
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636943256
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636943256
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636943256
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636943256
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp -25199
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_70
timestamp -25199
transform 1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_82
timestamp 1636943256
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_94
timestamp 1636943256
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_106
timestamp -25199
transform 1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_125
timestamp -25199
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_131
timestamp -25199
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_141
timestamp -25199
transform 1 0 14076 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636943256
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636943256
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636943256
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636943256
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636943256
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_65
timestamp -25199
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_71
timestamp -25199
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_75
timestamp -25199
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636943256
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1636943256
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1636943256
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp -25199
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp -25199
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp -25199
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636943256
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636943256
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636943256
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636943256
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636943256
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636943256
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636943256
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_93
timestamp -25199
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_99
timestamp -25199
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp -25199
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_122
timestamp -25199
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_130
timestamp -25199
transform 1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_142
timestamp -25199
transform 1 0 14168 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_148
timestamp -25199
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636943256
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636943256
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp -25199
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_35
timestamp -25199
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_66
timestamp 1636943256
transform 1 0 7176 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp -25199
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636943256
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp -25199
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_110
timestamp 1636943256
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_122
timestamp -25199
transform 1 0 12328 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp -25199
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636943256
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636943256
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636943256
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636943256
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp -25199
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp -25199
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_66
timestamp 1636943256
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_78
timestamp 1636943256
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_90
timestamp 1636943256
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp -25199
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp -25199
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636943256
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1636943256
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1636943256
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636943256
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636943256
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp -25199
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636943256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_41
timestamp -25199
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_70
timestamp 1636943256
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp -25199
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_99
timestamp 1636943256
transform 1 0 10212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_111
timestamp 1636943256
transform 1 0 11316 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_123
timestamp -25199
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp -25199
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp -25199
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636943256
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636943256
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636943256
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_39
timestamp -25199
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp -25199
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_67
timestamp -25199
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_91
timestamp -25199
transform 1 0 9476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp -25199
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636943256
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_125
timestamp -25199
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_148
timestamp -25199
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636943256
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636943256
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp -25199
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636943256
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636943256
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_53
timestamp -25199
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_61
timestamp 1636943256
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp -25199
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp -25199
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp -25199
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_108
timestamp 1636943256
transform 1 0 11040 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_120
timestamp -25199
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp -25199
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp -25199
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636943256
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636943256
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1636943256
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636943256
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp -25199
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp -25199
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636943256
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636943256
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636943256
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636943256
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp -25199
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp -25199
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636943256
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636943256
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1636943256
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636943256
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636943256
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1636943256
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_53
timestamp -25199
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_60
timestamp 1636943256
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_72
timestamp -25199
transform 1 0 7728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp -25199
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636943256
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636943256
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1636943256
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1636943256
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp -25199
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636943256
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636943256
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1636943256
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1636943256
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp -25199
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp -25199
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_66
timestamp 1636943256
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_78
timestamp 1636943256
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_90
timestamp 1636943256
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_102
timestamp -25199
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp -25199
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636943256
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636943256
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636943256
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636943256
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636943256
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp -25199
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636943256
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_41
timestamp -25199
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_45
timestamp -25199
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_71
timestamp -25199
transform 1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp -25199
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_93
timestamp -25199
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_114
timestamp -25199
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp -25199
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1636943256
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1636943256
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_39
timestamp -25199
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp -25199
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_71
timestamp -25199
transform 1 0 7636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_83
timestamp -25199
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_90
timestamp -25199
transform 1 0 9384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_94
timestamp -25199
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp -25199
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_117
timestamp -25199
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_142
timestamp -25199
transform 1 0 14168 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_148
timestamp -25199
transform 1 0 14720 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636943256
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636943256
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636943256
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_41
timestamp -25199
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_61
timestamp 1636943256
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_73
timestamp -25199
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp -25199
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_97
timestamp -25199
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_108
timestamp 1636943256
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_120
timestamp -25199
transform 1 0 12144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp -25199
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636943256
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636943256
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636943256
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1636943256
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp -25199
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp -25199
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1636943256
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1636943256
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1636943256
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1636943256
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp -25199
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp -25199
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636943256
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_125
timestamp -25199
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_142
timestamp -25199
transform 1 0 14168 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_148
timestamp -25199
transform 1 0 14720 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636943256
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636943256
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp -25199
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636943256
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1636943256
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_53
timestamp -25199
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_57
timestamp 1636943256
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_69
timestamp 1636943256
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp -25199
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636943256
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1636943256
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_109
timestamp -25199
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_113
timestamp 1636943256
transform 1 0 11500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_125
timestamp 1636943256
transform 1 0 12604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp -25199
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp -25199
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_25
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_26
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_27
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_28
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_29
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 15088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_30
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_31
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 15088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_32
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_33
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 15088 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_34
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_35
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_36
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_37
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_38
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_39
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 15088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_40
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 15088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_41
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 15088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_42
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_43
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_44
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_45
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_46
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 15088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_47
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_48
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 15088 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_49
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 15088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_53
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_55
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_56
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_70
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_71
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_72
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_73
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_74
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_76
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_78
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_79
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_80
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_81
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_82
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_83
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_84
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_85
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_86
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_87
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_88
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_89
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_90
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_91
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_92
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_93
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_94
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_95
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_96
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_97
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_98
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_100
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_101
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_103
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_104
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_105
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_106
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_107
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_108
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_109
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_110
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_111
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_112
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_113
timestamp -25199
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_114
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_115
timestamp -25199
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 15824 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 15824 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 15424 1368 16224 1488 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 15424 12928 16224 13048 0 FreeSans 480 0 0 0 clk_comp
port 3 nsew signal output
flabel metal3 s 15424 16328 16224 16448 0 FreeSans 480 0 0 0 clk_comp_shifted
port 4 nsew signal output
flabel metal3 s 15424 9528 16224 9648 0 FreeSans 480 0 0 0 dac_ctrl[0]
port 5 nsew signal output
flabel metal3 s 15424 7488 16224 7608 0 FreeSans 480 0 0 0 dac_ctrl[1]
port 6 nsew signal output
flabel metal3 s 15424 6808 16224 6928 0 FreeSans 480 0 0 0 dac_ctrl[2]
port 7 nsew signal output
flabel metal3 s 15424 13608 16224 13728 0 FreeSans 480 0 0 0 dac_ctrl[3]
port 8 nsew signal output
flabel metal3 s 15424 10208 16224 10328 0 FreeSans 480 0 0 0 dac_ctrl[4]
port 9 nsew signal output
flabel metal3 s 15424 5448 16224 5568 0 FreeSans 480 0 0 0 dac_ctrl[5]
port 10 nsew signal output
flabel metal3 s 15424 4768 16224 4888 0 FreeSans 480 0 0 0 dac_ctrl[6]
port 11 nsew signal output
flabel metal3 s 15424 8168 16224 8288 0 FreeSans 480 0 0 0 dac_ctrl[7]
port 12 nsew signal output
flabel metal3 s 15424 10888 16224 11008 0 FreeSans 480 0 0 0 dout[0]
port 13 nsew signal output
flabel metal3 s 15424 14288 16224 14408 0 FreeSans 480 0 0 0 dout[1]
port 14 nsew signal output
flabel metal3 s 15424 6128 16224 6248 0 FreeSans 480 0 0 0 dout[2]
port 15 nsew signal output
flabel metal3 s 15424 3408 16224 3528 0 FreeSans 480 0 0 0 dout[3]
port 16 nsew signal output
flabel metal3 s 15424 11568 16224 11688 0 FreeSans 480 0 0 0 dout[4]
port 17 nsew signal output
flabel metal3 s 15424 8848 16224 8968 0 FreeSans 480 0 0 0 dout[5]
port 18 nsew signal output
flabel metal3 s 15424 15648 16224 15768 0 FreeSans 480 0 0 0 dout[6]
port 19 nsew signal output
flabel metal3 s 15424 4088 16224 4208 0 FreeSans 480 0 0 0 dout[7]
port 20 nsew signal output
flabel metal3 s 15424 12248 16224 12368 0 FreeSans 480 0 0 0 en
port 21 nsew signal input
flabel metal3 s 15424 2728 16224 2848 0 FreeSans 480 0 0 0 samp
port 22 nsew signal output
flabel metal3 s 15424 2048 16224 2168 0 FreeSans 480 0 0 0 vcn
port 23 nsew signal input
flabel metal3 s 15424 14968 16224 15088 0 FreeSans 480 0 0 0 vcp
port 24 nsew signal input
rlabel metal1 8096 15232 8096 15232 0 VGND
rlabel metal1 8096 15776 8096 15776 0 VPWR
rlabel metal1 10212 13906 10212 13906 0 _000_
rlabel metal1 10442 10710 10442 10710 0 _001_
rlabel metal1 6210 12886 6210 12886 0 _002_
rlabel metal2 4738 9146 4738 9146 0 _003_
rlabel metal1 5888 13906 5888 13906 0 _004_
rlabel metal1 8464 10642 8464 10642 0 _005_
rlabel metal2 5750 10438 5750 10438 0 _006_
rlabel metal1 8924 13974 8924 13974 0 _007_
rlabel metal2 10442 8772 10442 8772 0 _008_
rlabel metal1 5934 6290 5934 6290 0 _009_
rlabel metal1 5888 6766 5888 6766 0 _010_
rlabel metal2 7774 6596 7774 6596 0 _011_
rlabel metal1 12880 10234 12880 10234 0 _012_
rlabel metal1 13340 13498 13340 13498 0 _013_
rlabel metal2 12742 6460 12742 6460 0 _014_
rlabel metal2 12466 13702 12466 13702 0 _015_
rlabel metal1 13110 10710 13110 10710 0 _016_
rlabel metal1 13340 8602 13340 8602 0 _017_
rlabel metal2 13202 14586 13202 14586 0 _018_
rlabel via1 13202 6717 13202 6717 0 _019_
rlabel metal1 11822 7412 11822 7412 0 _020_
rlabel metal1 12926 6698 12926 6698 0 _021_
rlabel metal1 4830 13838 4830 13838 0 _022_
rlabel metal1 11086 6426 11086 6426 0 _023_
rlabel metal1 7406 6732 7406 6732 0 _024_
rlabel metal2 9154 3468 9154 3468 0 _025_
rlabel metal1 10074 3502 10074 3502 0 _026_
rlabel metal2 8878 3502 8878 3502 0 _027_
rlabel metal1 9660 3502 9660 3502 0 _028_
rlabel metal1 12374 3570 12374 3570 0 _029_
rlabel metal1 13105 3502 13105 3502 0 _030_
rlabel via1 13289 3094 13289 3094 0 _031_
rlabel metal2 13478 13192 13478 13192 0 _032_
rlabel metal1 9246 3536 9246 3536 0 _033_
rlabel metal1 8464 6290 8464 6290 0 _034_
rlabel metal1 10810 10574 10810 10574 0 _035_
rlabel metal1 6992 13294 6992 13294 0 _036_
rlabel metal2 6670 12988 6670 12988 0 _037_
rlabel metal2 6854 9316 6854 9316 0 _038_
rlabel metal2 6578 9758 6578 9758 0 _039_
rlabel metal2 10534 6698 10534 6698 0 _040_
rlabel metal2 10350 6528 10350 6528 0 _041_
rlabel metal1 6394 13260 6394 13260 0 _042_
rlabel metal1 14030 12274 14030 12274 0 _043_
rlabel metal2 7038 13362 7038 13362 0 _044_
rlabel metal1 6900 12750 6900 12750 0 _045_
rlabel metal1 5750 13328 5750 13328 0 _046_
rlabel metal1 6854 6664 6854 6664 0 _047_
rlabel metal2 10074 10302 10074 10302 0 _048_
rlabel metal1 10488 10166 10488 10166 0 _049_
rlabel metal1 6808 9010 6808 9010 0 _050_
rlabel metal1 9476 13430 9476 13430 0 _051_
rlabel metal2 5474 13736 5474 13736 0 _052_
rlabel metal1 11224 6766 11224 6766 0 _053_
rlabel metal1 11270 13226 11270 13226 0 _054_
rlabel metal1 9982 13226 9982 13226 0 _055_
rlabel metal1 8556 10234 8556 10234 0 _056_
rlabel metal2 6762 10846 6762 10846 0 _057_
rlabel metal1 5934 10064 5934 10064 0 _058_
rlabel metal2 8418 13532 8418 13532 0 _059_
rlabel metal2 7130 9758 7130 9758 0 _060_
rlabel metal2 8694 13702 8694 13702 0 _061_
rlabel metal1 10626 8432 10626 8432 0 _062_
rlabel metal1 10902 8500 10902 8500 0 _063_
rlabel metal1 13662 13294 13662 13294 0 _064_
rlabel metal1 9246 3944 9246 3944 0 _065_
rlabel metal1 9154 3604 9154 3604 0 _066_
rlabel metal3 13946 1428 13946 1428 0 clk
rlabel metal2 13846 3910 13846 3910 0 clk_comp
rlabel metal2 12834 3604 12834 3604 0 clk_comp_shifted
rlabel metal2 11270 13498 11270 13498 0 cmp_processor_0.comp
rlabel via1 13100 10030 13100 10030 0 dac_ctrl[0]
rlabel metal1 13133 13294 13133 13294 0 dac_ctrl[1]
rlabel metal3 14084 6868 14084 6868 0 dac_ctrl[2]
rlabel via1 12640 13362 12640 13362 0 dac_ctrl[3]
rlabel metal1 14296 10574 14296 10574 0 dac_ctrl[4]
rlabel metal2 12374 6953 12374 6953 0 dac_ctrl[5]
rlabel metal1 11086 14586 11086 14586 0 dac_ctrl[6]
rlabel via1 13560 7378 13560 7378 0 dac_ctrl[7]
rlabel via2 13570 10965 13570 10965 0 dout[0]
rlabel metal2 14122 14195 14122 14195 0 dout[1]
rlabel via2 14122 6171 14122 6171 0 dout[2]
rlabel metal3 14268 3468 14268 3468 0 dout[3]
rlabel metal2 14582 11169 14582 11169 0 dout[4]
rlabel metal2 13938 8857 13938 8857 0 dout[5]
rlabel metal2 14030 15385 14030 15385 0 dout[6]
rlabel metal3 14728 4148 14728 4148 0 dout[7]
rlabel metal1 13202 4046 13202 4046 0 en
rlabel via2 9890 2805 9890 2805 0 samp
rlabel metal1 7912 13294 7912 13294 0 sar_logic_0.count\[0\]
rlabel metal1 6762 13430 6762 13430 0 sar_logic_0.count\[1\]
rlabel metal2 6486 13600 6486 13600 0 sar_logic_0.count\[2\]
rlabel metal1 7452 13226 7452 13226 0 sar_logic_0.eoc
rlabel metal1 10856 4658 10856 4658 0 smp_clk_div_0.start
rlabel metal1 14030 3502 14030 3502 0 vcn
rlabel metal2 13938 13617 13938 13617 0 vcp
<< properties >>
string FIXED_BBOX 0 0 20000 40000
<< end >>
