magic
tech sky130A
magscale 1 2
timestamp 1722275549
use sky130_fd_pr__nfet_01v8_QJTADH  sky130_fd_pr__nfet_01v8_QJTADH_0
timestamp 1722275450
transform 1 0 1612 0 1 -393
box -558 -167 558 167
use sky130_fd_pr__nfet_01v8_QJTADH  sky130_fd_pr__nfet_01v8_QJTADH_1
timestamp 1722275450
transform -1 0 1614 0 -1 -795
box -558 -167 558 167
use sky130_fd_pr__pfet_01v8_XEBJEJ  sky130_fd_pr__pfet_01v8_XEBJEJ_0
timestamp 1722275450
transform 1 0 1112 0 1 122
box -1094 -264 1094 298
use sky130_fd_pr__pfet_01v8_XEBJEJ  sky130_fd_pr__pfet_01v8_XEBJEJ_1
timestamp 1722275450
transform -1 0 1112 0 -1 986
box -1094 -264 1094 298
<< end >>
